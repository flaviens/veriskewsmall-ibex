// Copyright lowRISC contributors.
// Copyright 2017 ETH Zurich and University of Bologna, see also CREDITS.md.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

/**
 * Package with constants used by Ibex
 */
package ibex_pkg;

////////////////
// IO Structs //
////////////////

typedef struct packed {
  logic [31:0] current_pc;
  logic [31:0] next_pc;
  logic [31:0] last_data_addr;
  logic [31:0] exception_addr;
} crash_dump_t;

typedef struct packed {
  logic        dummy_instr_id;
  logic [4:0]  raddr_a;
  logic [4:0]  waddr_a;
  logic        we_a;
  logic [4:0]  raddr_b;
} core2rf_t;

/////////////////////
// Parameter Enums //
/////////////////////

typedef enum integer {
  RegFileFF    = 0,
  RegFileFPGA  = 1,
  RegFileLatch = 2
} regfile_e;

typedef enum integer {
  RV32MNone        = 0,
  RV32MSlow        = 1,
  RV32MFast        = 2,
  RV32MSingleCycle = 3
} rv32m_e;

typedef enum integer {
  RV32BNone     = 0,
  RV32BBalanced = 1,
  RV32BFull     = 2
} rv32b_e;

/////////////
// Opcodes //
/////////////

typedef enum logic [6:0] {
  OPCODE_LOAD     = 7'h03,
  OPCODE_MISC_MEM = 7'h0f,
  OPCODE_OP_IMM   = 7'h13,
  OPCODE_AUIPC    = 7'h17,
  OPCODE_STORE    = 7'h23,
  OPCODE_OP       = 7'h33,
  OPCODE_LUI      = 7'h37,
  OPCODE_BRANCH   = 7'h63,
  OPCODE_JALR     = 7'h67,
  OPCODE_JAL      = 7'h6f,
  OPCODE_SYSTEM   = 7'h73
} opcode_e;


////////////////////
// ALU operations //
////////////////////

typedef enum logic [5:0] {
  // Arithmetics
  ALU_ADD,
  ALU_SUB,

  // Logics
  ALU_XOR,
  ALU_OR,
  ALU_AND,
  // RV32B
  ALU_XNOR,
  ALU_ORN,
  ALU_ANDN,

  // Shifts
  ALU_SRA,
  ALU_SRL,
  ALU_SLL,
  // RV32B
  ALU_SRO,
  ALU_SLO,
  ALU_ROR,
  ALU_ROL,
  ALU_GREV,
  ALU_GORC,
  ALU_SHFL,
  ALU_UNSHFL,

  // Comparisons
  ALU_LT,
  ALU_LTU,
  ALU_GE,
  ALU_GEU,
  ALU_EQ,
  ALU_NE,
  // RV32B
  ALU_MIN,
  ALU_MINU,
  ALU_MAX,
  ALU_MAXU,

  // Pack
  // RV32B
  ALU_PACK,
  ALU_PACKU,
  ALU_PACKH,

  // Sign-Extend
  // RV32B
  ALU_SEXTB,
  ALU_SEXTH,

  // Bitcounting
  // RV32B
  ALU_CLZ,
  ALU_CTZ,
  ALU_PCNT,

  // Set lower than
  ALU_SLT,
  ALU_SLTU,

  // Ternary Bitmanip Operations
  // RV32B
  ALU_CMOV,
  ALU_CMIX,
  ALU_FSL,
  ALU_FSR,

  // Single-Bit Operations
  // RV32B
  ALU_SBSET,
  ALU_SBCLR,
  ALU_SBINV,
  ALU_SBEXT,

  // Bit Extract / Deposit
  // RV32B
  ALU_BEXT,
  ALU_BDEP,

  // Bit Field Place
  // RV32B
  ALU_BFP,

  // Carry-less Multiply
  // RV32B
  ALU_CLMUL,
  ALU_CLMULR,
  ALU_CLMULH,

  // Cyclic Redundancy Check
  ALU_CRC32_B,
  ALU_CRC32C_B,
  ALU_CRC32_H,
  ALU_CRC32C_H,
  ALU_CRC32_W,
  ALU_CRC32C_W
} alu_op_e;

typedef enum logic [1:0] {
  // Multiplier/divider
  MD_OP_MULL,
  MD_OP_MULH,
  MD_OP_DIV,
  MD_OP_REM
} md_op_e;


//////////////////////////////////
// Control and status registers //
//////////////////////////////////

// CSR operations
typedef enum logic [1:0] {
  CSR_OP_READ,
  CSR_OP_WRITE,
  CSR_OP_SET,
  CSR_OP_CLEAR
} csr_op_e;

// Privileged mode
typedef enum logic[1:0] {
  PRIV_LVL_M = 2'b11,
  PRIV_LVL_H = 2'b10,
  PRIV_LVL_S = 2'b01,
  PRIV_LVL_U = 2'b00
} priv_lvl_e;

// Constants for the dcsr.xdebugver fields
typedef enum logic[3:0] {
   XDEBUGVER_NO     = 4'd0, // no external debug support
   XDEBUGVER_STD    = 4'd4, // external debug according to RISC-V debug spec
   XDEBUGVER_NONSTD = 4'd15 // debug not conforming to RISC-V debug spec
} x_debug_ver_e;

//////////////
// WB stage //
//////////////

// Type of instruction present in writeback stage
typedef enum logic[1:0] {
  WB_INSTR_LOAD,  // Instruction is awaiting load data
  WB_INSTR_STORE, // Instruction is awaiting store response
  WB_INSTR_OTHER  // Instruction doesn't fit into above categories
} wb_instr_type_e;

//////////////
// ID stage //
//////////////

// Operand a selection
typedef enum logic[1:0] {
  OP_A_REG_A,
  OP_A_FWD,
  OP_A_CURRPC,
  OP_A_IMM
} op_a_sel_e;

// Immediate a selection
typedef enum logic {
  IMM_A_Z,
  IMM_A_ZERO
} imm_a_sel_e;

// Operand b selection
typedef enum logic {
  OP_B_REG_B,
  OP_B_IMM
} op_b_sel_e;

// Immediate b selection
typedef enum logic [2:0] {
  IMM_B_I,
  IMM_B_S,
  IMM_B_B,
  IMM_B_U,
  IMM_B_J,
  IMM_B_INCR_PC,
  IMM_B_INCR_ADDR
} imm_b_sel_e;

// Regfile write data selection
typedef enum logic {
  RF_WD_EX,
  RF_WD_CSR
} rf_wd_sel_e;

//////////////
// IF stage //
//////////////

// PC mux selection
typedef enum logic [2:0] {
  PC_BOOT,
  PC_JUMP,
  PC_EXC,
  PC_ERET,
  PC_DRET,
  PC_BP
} pc_sel_e;

// Exception PC mux selection
typedef enum logic [1:0] {
  EXC_PC_EXC,
  EXC_PC_IRQ,
  EXC_PC_DBD,
  EXC_PC_DBG_EXC // Exception while in debug mode
} exc_pc_sel_e;

// Interrupt requests
typedef struct packed {
  logic        irq_software;
  logic        irq_timer;
  logic        irq_external;
  logic [14:0] irq_fast; // 15 fast interrupts,
                         // one interrupt is reserved for NMI (not visible through mip/mie)
} irqs_t;

// Exception cause
typedef enum logic [5:0] {
  EXC_CAUSE_IRQ_SOFTWARE_M     = {1'b1, 5'd03},
  EXC_CAUSE_IRQ_TIMER_M        = {1'b1, 5'd07},
  EXC_CAUSE_IRQ_EXTERNAL_M     = {1'b1, 5'd11},
  // EXC_CAUSE_IRQ_FAST_0      = {1'b1, 5'd16},
  // EXC_CAUSE_IRQ_FAST_14     = {1'b1, 5'd30},
  EXC_CAUSE_IRQ_NM             = {1'b1, 5'd31}, // == EXC_CAUSE_IRQ_FAST_15
  EXC_CAUSE_INSN_ADDR_MISA     = {1'b0, 5'd00},
  EXC_CAUSE_INSTR_ACCESS_FAULT = {1'b0, 5'd01},
  EXC_CAUSE_ILLEGAL_INSN       = {1'b0, 5'd02},
  EXC_CAUSE_BREAKPOINT         = {1'b0, 5'd03},
  EXC_CAUSE_LOAD_ACCESS_FAULT  = {1'b0, 5'd05},
  EXC_CAUSE_STORE_ACCESS_FAULT = {1'b0, 5'd07},
  EXC_CAUSE_ECALL_UMODE        = {1'b0, 5'd08},
  EXC_CAUSE_ECALL_MMODE        = {1'b0, 5'd11}
} exc_cause_e;

// Debug cause
typedef enum logic [2:0] {
  DBG_CAUSE_NONE    = 3'h0,
  DBG_CAUSE_EBREAK  = 3'h1,
  DBG_CAUSE_TRIGGER = 3'h2,
  DBG_CAUSE_HALTREQ = 3'h3,
  DBG_CAUSE_STEP    = 3'h4
} dbg_cause_e;

// ICache constants
parameter int unsigned ADDR_W          = 32;
parameter int unsigned BUS_SIZE        = 32;
parameter int unsigned BUS_BYTES       = BUS_SIZE/8;
parameter int unsigned BUS_W           = $clog2(BUS_BYTES);
parameter int unsigned IC_SIZE_BYTES   = 4096;
parameter int unsigned IC_NUM_WAYS     = 2;
parameter int unsigned IC_LINE_SIZE    = 64;
parameter int unsigned IC_LINE_BYTES   = IC_LINE_SIZE/8;
parameter int unsigned IC_LINE_W       = $clog2(IC_LINE_BYTES);
parameter int unsigned IC_NUM_LINES    = IC_SIZE_BYTES / IC_NUM_WAYS / IC_LINE_BYTES;
parameter int unsigned IC_LINE_BEATS   = IC_LINE_BYTES / BUS_BYTES;
parameter int unsigned IC_LINE_BEATS_W = $clog2(IC_LINE_BEATS);
parameter int unsigned IC_INDEX_W      = $clog2(IC_NUM_LINES);
parameter int unsigned IC_INDEX_HI     = IC_INDEX_W + IC_LINE_W - 1;
parameter int unsigned IC_TAG_SIZE     = ADDR_W - IC_INDEX_W - IC_LINE_W + 1; // 1 valid bit
parameter int unsigned IC_OUTPUT_BEATS = (BUS_BYTES / 2); // number of halfwords

// PMP constants
parameter int unsigned PMP_MAX_REGIONS      = 16;
parameter int unsigned PMP_CFG_W            = 8;

// PMP acces type
parameter int unsigned PMP_I = 0;
parameter int unsigned PMP_D = 1;

typedef enum logic [1:0] {
  PMP_ACC_EXEC    = 2'b00,
  PMP_ACC_WRITE   = 2'b01,
  PMP_ACC_READ    = 2'b10
} pmp_req_e;

// PMP cfg structures
typedef enum logic [1:0] {
  PMP_MODE_OFF   = 2'b00,
  PMP_MODE_TOR   = 2'b01,
  PMP_MODE_NA4   = 2'b10,
  PMP_MODE_NAPOT = 2'b11
} pmp_cfg_mode_e;

typedef struct packed {
  logic          lock;
  pmp_cfg_mode_e mode;
  logic          exec;
  logic          write;
  logic          read;
} pmp_cfg_t;

// Machine Security Configuration (ePMP)
typedef struct packed {
  logic rlb;  // Rule Locking Bypass
  logic mmwp; // Machine Mode Whitelist Policy
  logic mml;  // Machine Mode Lockdown
} pmp_mseccfg_t;

// CSRs
typedef enum logic[11:0] {
  // Machine information
  CSR_MHARTID   = 12'hF14,

  // Machine trap setup
  CSR_MSTATUS   = 12'h300,
  CSR_MISA      = 12'h301,
  CSR_MIE       = 12'h304,
  CSR_MTVEC     = 12'h305,
  CSR_MCOUNTEREN= 12'h306,

  // Machine trap handling
  CSR_MSCRATCH  = 12'h340,
  CSR_MEPC      = 12'h341,
  CSR_MCAUSE    = 12'h342,
  CSR_MTVAL     = 12'h343,
  CSR_MIP       = 12'h344,

  CSR_MSECCFG   = 12'h390,
  CSR_MSECCFGH  = 12'h391,

  // Physical memory protection
  CSR_PMPCFG0   = 12'h3A0,
  CSR_PMPCFG1   = 12'h3A1,
  CSR_PMPCFG2   = 12'h3A2,
  CSR_PMPCFG3   = 12'h3A3,
  CSR_PMPADDR0  = 12'h3B0,
  CSR_PMPADDR1  = 12'h3B1,
  CSR_PMPADDR2  = 12'h3B2,
  CSR_PMPADDR3  = 12'h3B3,
  CSR_PMPADDR4  = 12'h3B4,
  CSR_PMPADDR5  = 12'h3B5,
  CSR_PMPADDR6  = 12'h3B6,
  CSR_PMPADDR7  = 12'h3B7,
  CSR_PMPADDR8  = 12'h3B8,
  CSR_PMPADDR9  = 12'h3B9,
  CSR_PMPADDR10 = 12'h3BA,
  CSR_PMPADDR11 = 12'h3BB,
  CSR_PMPADDR12 = 12'h3BC,
  CSR_PMPADDR13 = 12'h3BD,
  CSR_PMPADDR14 = 12'h3BE,
  CSR_PMPADDR15 = 12'h3BF,

  // Debug trigger
  CSR_TSELECT   = 12'h7A0,
  CSR_TDATA1    = 12'h7A1,
  CSR_TDATA2    = 12'h7A2,
  CSR_TDATA3    = 12'h7A3,
  CSR_MCONTEXT  = 12'h7A8,
  CSR_SCONTEXT  = 12'h7AA,

  // Debug/trace
  CSR_DCSR      = 12'h7b0,
  CSR_DPC       = 12'h7b1,

  // Debug
  CSR_DSCRATCH0 = 12'h7b2, // optional
  CSR_DSCRATCH1 = 12'h7b3, // optional

  // Machine Counter/Timers
  CSR_MCOUNTINHIBIT  = 12'h320,
  CSR_MHPMEVENT3     = 12'h323,
  CSR_MHPMEVENT4     = 12'h324,
  CSR_MHPMEVENT5     = 12'h325,
  CSR_MHPMEVENT6     = 12'h326,
  CSR_MHPMEVENT7     = 12'h327,
  CSR_MHPMEVENT8     = 12'h328,
  CSR_MHPMEVENT9     = 12'h329,
  CSR_MHPMEVENT10    = 12'h32A,
  CSR_MHPMEVENT11    = 12'h32B,
  CSR_MHPMEVENT12    = 12'h32C,
  CSR_MHPMEVENT13    = 12'h32D,
  CSR_MHPMEVENT14    = 12'h32E,
  CSR_MHPMEVENT15    = 12'h32F,
  CSR_MHPMEVENT16    = 12'h330,
  CSR_MHPMEVENT17    = 12'h331,
  CSR_MHPMEVENT18    = 12'h332,
  CSR_MHPMEVENT19    = 12'h333,
  CSR_MHPMEVENT20    = 12'h334,
  CSR_MHPMEVENT21    = 12'h335,
  CSR_MHPMEVENT22    = 12'h336,
  CSR_MHPMEVENT23    = 12'h337,
  CSR_MHPMEVENT24    = 12'h338,
  CSR_MHPMEVENT25    = 12'h339,
  CSR_MHPMEVENT26    = 12'h33A,
  CSR_MHPMEVENT27    = 12'h33B,
  CSR_MHPMEVENT28    = 12'h33C,
  CSR_MHPMEVENT29    = 12'h33D,
  CSR_MHPMEVENT30    = 12'h33E,
  CSR_MHPMEVENT31    = 12'h33F,
  CSR_MCYCLE         = 12'hB00,
  CSR_MINSTRET       = 12'hB02,
  CSR_MHPMCOUNTER3   = 12'hB03,
  CSR_MHPMCOUNTER4   = 12'hB04,
  CSR_MHPMCOUNTER5   = 12'hB05,
  CSR_MHPMCOUNTER6   = 12'hB06,
  CSR_MHPMCOUNTER7   = 12'hB07,
  CSR_MHPMCOUNTER8   = 12'hB08,
  CSR_MHPMCOUNTER9   = 12'hB09,
  CSR_MHPMCOUNTER10  = 12'hB0A,
  CSR_MHPMCOUNTER11  = 12'hB0B,
  CSR_MHPMCOUNTER12  = 12'hB0C,
  CSR_MHPMCOUNTER13  = 12'hB0D,
  CSR_MHPMCOUNTER14  = 12'hB0E,
  CSR_MHPMCOUNTER15  = 12'hB0F,
  CSR_MHPMCOUNTER16  = 12'hB10,
  CSR_MHPMCOUNTER17  = 12'hB11,
  CSR_MHPMCOUNTER18  = 12'hB12,
  CSR_MHPMCOUNTER19  = 12'hB13,
  CSR_MHPMCOUNTER20  = 12'hB14,
  CSR_MHPMCOUNTER21  = 12'hB15,
  CSR_MHPMCOUNTER22  = 12'hB16,
  CSR_MHPMCOUNTER23  = 12'hB17,
  CSR_MHPMCOUNTER24  = 12'hB18,
  CSR_MHPMCOUNTER25  = 12'hB19,
  CSR_MHPMCOUNTER26  = 12'hB1A,
  CSR_MHPMCOUNTER27  = 12'hB1B,
  CSR_MHPMCOUNTER28  = 12'hB1C,
  CSR_MHPMCOUNTER29  = 12'hB1D,
  CSR_MHPMCOUNTER30  = 12'hB1E,
  CSR_MHPMCOUNTER31  = 12'hB1F,
  CSR_MCYCLEH        = 12'hB80,
  CSR_MINSTRETH      = 12'hB82,
  CSR_MHPMCOUNTER3H  = 12'hB83,
  CSR_MHPMCOUNTER4H  = 12'hB84,
  CSR_MHPMCOUNTER5H  = 12'hB85,
  CSR_MHPMCOUNTER6H  = 12'hB86,
  CSR_MHPMCOUNTER7H  = 12'hB87,
  CSR_MHPMCOUNTER8H  = 12'hB88,
  CSR_MHPMCOUNTER9H  = 12'hB89,
  CSR_MHPMCOUNTER10H = 12'hB8A,
  CSR_MHPMCOUNTER11H = 12'hB8B,
  CSR_MHPMCOUNTER12H = 12'hB8C,
  CSR_MHPMCOUNTER13H = 12'hB8D,
  CSR_MHPMCOUNTER14H = 12'hB8E,
  CSR_MHPMCOUNTER15H = 12'hB8F,
  CSR_MHPMCOUNTER16H = 12'hB90,
  CSR_MHPMCOUNTER17H = 12'hB91,
  CSR_MHPMCOUNTER18H = 12'hB92,
  CSR_MHPMCOUNTER19H = 12'hB93,
  CSR_MHPMCOUNTER20H = 12'hB94,
  CSR_MHPMCOUNTER21H = 12'hB95,
  CSR_MHPMCOUNTER22H = 12'hB96,
  CSR_MHPMCOUNTER23H = 12'hB97,
  CSR_MHPMCOUNTER24H = 12'hB98,
  CSR_MHPMCOUNTER25H = 12'hB99,
  CSR_MHPMCOUNTER26H = 12'hB9A,
  CSR_MHPMCOUNTER27H = 12'hB9B,
  CSR_MHPMCOUNTER28H = 12'hB9C,
  CSR_MHPMCOUNTER29H = 12'hB9D,
  CSR_MHPMCOUNTER30H = 12'hB9E,
  CSR_MHPMCOUNTER31H = 12'hB9F,
  CSR_CPUCTRL        = 12'h7C0,
  CSR_SECURESEED     = 12'h7C1
} csr_num_e;

// CSR pmp-related offsets
parameter logic [11:0] CSR_OFF_PMP_CFG  = 12'h3A0; // pmp_cfg  @ 12'h3a0 - 12'h3a3
parameter logic [11:0] CSR_OFF_PMP_ADDR = 12'h3B0; // pmp_addr @ 12'h3b0 - 12'h3bf

// CSR status bits
parameter int unsigned CSR_MSTATUS_MIE_BIT      = 3;
parameter int unsigned CSR_MSTATUS_MPIE_BIT     = 7;
parameter int unsigned CSR_MSTATUS_MPP_BIT_LOW  = 11;
parameter int unsigned CSR_MSTATUS_MPP_BIT_HIGH = 12;
parameter int unsigned CSR_MSTATUS_MPRV_BIT     = 17;
parameter int unsigned CSR_MSTATUS_TW_BIT       = 21;

// CSR machine ISA
parameter logic [1:0] CSR_MISA_MXL = 2'd1; // M-XLEN: XLEN in M-Mode for RV32

// CSR interrupt pending/enable bits
parameter int unsigned CSR_MSIX_BIT      = 3;
parameter int unsigned CSR_MTIX_BIT      = 7;
parameter int unsigned CSR_MEIX_BIT      = 11;
parameter int unsigned CSR_MFIX_BIT_LOW  = 16;
parameter int unsigned CSR_MFIX_BIT_HIGH = 30;

// CSR Machine Security Configuration bits
parameter int unsigned CSR_MSECCFG_MML_BIT  = 0;
parameter int unsigned CSR_MSECCFG_MMWP_BIT = 1;
parameter int unsigned CSR_MSECCFG_RLB_BIT  = 2;

endpackage


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0


/**
 * Utility functions
 */
package prim_util_pkg;
  /**
   * Math function: $clog2 as specified in Verilog-2005
   *
   * Do not use this function if $clog2() is available.
   *
   * clog2 =          0        for value == 0
   *         ceil(log2(value)) for value >= 1
   *
   * This implementation is a synthesizable variant of the $clog2 function as
   * specified in the Verilog-2005 standard (IEEE 1364-2005).
   *
   * To quote the standard:
   *   The system function $clog2 shall return the ceiling of the log
   *   base 2 of the argument (the log rounded up to an integer
   *   value). The argument can be an integer or an arbitrary sized
   *   vector value. The argument shall be treated as an unsigned
   *   value, and an argument value of 0 shall produce a result of 0.
   */
  function automatic integer _clog2(integer value);
    integer result;
    // Use an intermediate value to avoid assigning to an input port, which produces a warning in
    // Synopsys DC.
    integer v = value;
    v = v - 1;
    for (result = 0; v > 0; result++) begin
      v = v >> 1;
    end
    return result;
  endfunction


  /**
   * Math function: Number of bits needed to address |value| items.
   *
   *                  0        for value == 0
   * vbits =          1        for value == 1
   *         ceil(log2(value)) for value > 1
   *
   *
   * The primary use case for this function is the definition of registers/arrays
   * which are wide enough to contain |value| items.
   *
   * This function identical to $clog2() for all input values except the value 1;
   * it could be considered an "enhanced" $clog2() function.
   *
   *
   * Example 1:
   *   parameter Items = 1;
   *   localparam ItemsWidth = vbits(Items); // 1
   *   logic [ItemsWidth-1:0] item_register; // items_register is now [0:0]
   *
   * Example 2:
   *   parameter Items = 64;
   *   localparam ItemsWidth = vbits(Items); // 6
   *   logic [ItemsWidth-1:0] item_register; // items_register is now [5:0]
   *
   * Note: If you want to store the number "value" inside a register, you need
   * a register with size vbits(value + 1), since you also need to store
   * the number 0.
   *
   * Example 3:
   *   logic [vbits(64)-1:0]     store_64_logic_values; // width is [5:0]
   *   logic [vbits(64 + 1)-1:0] store_number_64;       // width is [6:0]
   */
  function automatic integer vbits(integer value);
`ifdef XCELIUM
    // The use of system functions was not allowed here in Verilog-2001, but is
    // valid since (System)Verilog-2005, which is also when $clog2() first
    // appeared.
    // Xcelium < 19.10 does not yet support the use of $clog2() here, fall back
    // to an implementation without a system function. Remove this workaround
    // if we require a newer Xcelium version.
    // See #2579 and #2597.
    return (value == 1) ? 1 : _clog2(value);
`else
    return (value == 1) ? 1 : $clog2(value);
`endif
  endfunction

endpackage

// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Life cycle state encoding definition.
//
// DO NOT EDIT THIS FILE DIRECTLY.
// It has been generated with
// $ ./util/design/gen-lc-state-enc.py --seed 10167336684108184581
//
package lc_ctrl_state_pkg;

  import prim_util_pkg::vbits;

  ///////////////////////////////
  // General size declarations //
  ///////////////////////////////

  parameter int LcValueWidth = 16;

  parameter int NumLcStateValues = 12;
  parameter int LcStateWidth = NumLcStateValues * LcValueWidth;
  parameter int NumLcStates = 13;
  parameter int DecLcStateWidth = vbits(NumLcStates);

  parameter int NumLcCountValues = 16;
  parameter int LcCountWidth = NumLcCountValues * LcValueWidth;
  parameter int NumLcCountStates = 17;
  parameter int DecLcCountWidth = vbits(NumLcCountStates);

  parameter int NumLcIdStateValues = 1;
  parameter int LcIdStateWidth = NumLcIdStateValues * LcValueWidth;
  parameter int NumLcIdStates = 2;
  parameter int DecLcIdStateWidth = vbits(NumLcIdStates+1);

  /////////////////////////////////////////////
  // Life cycle manufacturing state encoding //
  /////////////////////////////////////////////

  // These values have been generated such that they are incrementally writeable with respect
  // to the ECC polynomial specified. The values are used to define the life cycle manufacturing
  // state and transition counter encoding in lc_ctrl_pkg.sv.
  //
  // The values are unique and have the following statistics (considering all 16
  // data and 6 ECC bits):
  //
  // - Minimum Hamming weight: 8
  // - Maximum Hamming weight: 16
  // - Minimum Hamming distance from any other value: 6
  // - Maximum Hamming distance from any other value: 20
  //
  // Hamming distance histogram:
  //
  //  0: --
  //  1: --
  //  2: --
  //  3: --
  //  4: --
  //  5: --
  //  6: |||| (6.84%)
  //  7: --
  //  8: ||||||||||| (16.70%)
  //  9: --
  // 10: ||||||||||||||||||| (29.10%)
  // 11: --
  // 12: |||||||||||||||||||| (29.82%)
  // 13: --
  // 14: |||||||| (12.83%)
  // 15: --
  // 16: || (4.30%)
  // 17: --
  // 18:  (0.36%)
  // 19: --
  // 20:  (0.06%)
  // 21: --
  // 22: --
  //
  //
  // Note that the ECC bits are not defined in this package as they will be calculated by
  // the OTP ECC logic at runtime.

  // The A/B values are used for the encoded LC state.
  parameter logic [15:0] A0 = 16'b1000011000111000; // ECC: 6'b110000
  parameter logic [15:0] B0 = 16'b1110011001111001; // ECC: 6'b111111

  parameter logic [15:0] A1 = 16'b1100011000100110; // ECC: 6'b101001
  parameter logic [15:0] B1 = 16'b1101111101101110; // ECC: 6'b101011

  parameter logic [15:0] A2 = 16'b0010000111101100; // ECC: 6'b110010
  parameter logic [15:0] B2 = 16'b0111011111101101; // ECC: 6'b110110

  parameter logic [15:0] A3 = 16'b0001100111101000; // ECC: 6'b000100
  parameter logic [15:0] B3 = 16'b1101101111101100; // ECC: 6'b001101

  parameter logic [15:0] A4 = 16'b1001011001100100; // ECC: 6'b000001
  parameter logic [15:0] B4 = 16'b1101111001110100; // ECC: 6'b101101

  parameter logic [15:0] A5 = 16'b0001011000010110; // ECC: 6'b111001
  parameter logic [15:0] B5 = 16'b1011011001110111; // ECC: 6'b111101

  parameter logic [15:0] A6 = 16'b0101001001010010; // ECC: 6'b001111
  parameter logic [15:0] B6 = 16'b1101111111110010; // ECC: 6'b001111

  parameter logic [15:0] A7 = 16'b0010001001011111; // ECC: 6'b011000
  parameter logic [15:0] B7 = 16'b0011101011111111; // ECC: 6'b011101

  parameter logic [15:0] A8 = 16'b0000001110111001; // ECC: 6'b001000
  parameter logic [15:0] B8 = 16'b1100001110111111; // ECC: 6'b101010

  parameter logic [15:0] A9 = 16'b1100100101111000; // ECC: 6'b010010
  parameter logic [15:0] B9 = 16'b1111101101111001; // ECC: 6'b011110

  parameter logic [15:0] A10 = 16'b0010000110110111; // ECC: 6'b010001
  parameter logic [15:0] B10 = 16'b1011010111111111; // ECC: 6'b010101

  parameter logic [15:0] A11 = 16'b1011000100000111; // ECC: 6'b011001
  parameter logic [15:0] B11 = 16'b1111110110000111; // ECC: 6'b011111


  // The C/D values are used for the encoded LC transition counter.
  parameter logic [15:0] C0 = 16'b0011100000010000; // ECC: 6'b111001
  parameter logic [15:0] D0 = 16'b1111100100110000; // ECC: 6'b111111

  parameter logic [15:0] C1 = 16'b0011000010101011; // ECC: 6'b100110
  parameter logic [15:0] D1 = 16'b1011010011111011; // ECC: 6'b111110

  parameter logic [15:0] C2 = 16'b0011110100100000; // ECC: 6'b011000
  parameter logic [15:0] D2 = 16'b0011111101101011; // ECC: 6'b011100

  parameter logic [15:0] C3 = 16'b1010101100010010; // ECC: 6'b111000
  parameter logic [15:0] D3 = 16'b1111111110011010; // ECC: 6'b111010

  parameter logic [15:0] C4 = 16'b0100011010010100; // ECC: 6'b110110
  parameter logic [15:0] D4 = 16'b0101111110010111; // ECC: 6'b111110

  parameter logic [15:0] C5 = 16'b1011111110000101; // ECC: 6'b000000
  parameter logic [15:0] D5 = 16'b1011111111010111; // ECC: 6'b000111

  parameter logic [15:0] C6 = 16'b1110010000010111; // ECC: 6'b010100
  parameter logic [15:0] D6 = 16'b1111110010111111; // ECC: 6'b010110

  parameter logic [15:0] C7 = 16'b0100100101011010; // ECC: 6'b001000
  parameter logic [15:0] D7 = 16'b1110100111111111; // ECC: 6'b001101

  parameter logic [15:0] C8 = 16'b0000110000011011; // ECC: 6'b110110
  parameter logic [15:0] D8 = 16'b0011111000011111; // ECC: 6'b111111

  parameter logic [15:0] C9 = 16'b0111001100010100; // ECC: 6'b011001
  parameter logic [15:0] D9 = 16'b1111101101110110; // ECC: 6'b111001

  parameter logic [15:0] C10 = 16'b0001101110100010; // ECC: 6'b100011
  parameter logic [15:0] D10 = 16'b0011111111100011; // ECC: 6'b110111

  parameter logic [15:0] C11 = 16'b0000110101000010; // ECC: 6'b111101
  parameter logic [15:0] D11 = 16'b1100110111010110; // ECC: 6'b111111

  parameter logic [15:0] C12 = 16'b0001111111010001; // ECC: 6'b000010
  parameter logic [15:0] D12 = 16'b0001111111111001; // ECC: 6'b101111

  parameter logic [15:0] C13 = 16'b0010010000110000; // ECC: 6'b111111
  parameter logic [15:0] D13 = 16'b0111011100110101; // ECC: 6'b111111

  parameter logic [15:0] C14 = 16'b0010111010001111; // ECC: 6'b001000
  parameter logic [15:0] D14 = 16'b1011111010111111; // ECC: 6'b101100

  parameter logic [15:0] C15 = 16'b0100010000111101; // ECC: 6'b011010
  parameter logic [15:0] D15 = 16'b0101110011111101; // ECC: 6'b111110


  // The E/F values are used for the encoded ID state.
  parameter logic [15:0] E0 = 16'b1110000000101100; // ECC: 6'b111001
  parameter logic [15:0] F0 = 16'b1110010110111101; // ECC: 6'b111101


  parameter logic [15:0] ZRO = 16'h0;

  ////////////////////////
  // Derived enum types //
  ////////////////////////

  typedef enum logic [LcStateWidth-1:0] {
    LcStRaw           = {ZRO, ZRO, ZRO, ZRO, ZRO, ZRO, ZRO, ZRO, ZRO, ZRO, ZRO, ZRO},
    LcStTestUnlocked0 = {A11, A10,  A9,  A8,  A7,  A6,  A5,  A4,  A3,  A2,  A1,  B0},
    LcStTestLocked0   = {A11, A10,  A9,  A8,  A7,  A6,  A5,  A4,  A3,  A2,  B1,  B0},
    LcStTestUnlocked1 = {A11, A10,  A9,  A8,  A7,  A6,  A5,  A4,  A3,  B2,  B1,  B0},
    LcStTestLocked1   = {A11, A10,  A9,  A8,  A7,  A6,  A5,  A4,  B3,  B2,  B1,  B0},
    LcStTestUnlocked2 = {A11, A10,  A9,  A8,  A7,  A6,  A5,  B4,  B3,  B2,  B1,  B0},
    LcStTestLocked2   = {A11, A10,  A9,  A8,  A7,  A6,  B5,  B4,  B3,  B2,  B1,  B0},
    LcStTestUnlocked3 = {A11, A10,  A9,  A8,  A7,  B6,  B5,  B4,  B3,  B2,  B1,  B0},
    LcStDev           = {A11, A10,  A9,  A8,  B7,  B6,  B5,  B4,  B3,  B2,  B1,  B0},
    LcStProd          = {A11, A10,  A9,  B8,  A7,  B6,  B5,  B4,  B3,  B2,  B1,  B0},
    LcStProdEnd       = {A11, A10,  B9,  A8,  A7,  B6,  B5,  B4,  B3,  B2,  B1,  B0},
    LcStRma           = {B11, B10,  A9,  B8,  B7,  B6,  B5,  B4,  B3,  B2,  B1,  B0},
    LcStScrap         = {B11, B10,  B9,  B8,  B7,  B6,  B5,  B4,  B3,  B2,  B1,  B0}
  } lc_state_e;

  typedef enum logic [LcIdStateWidth-1:0] {
    LcIdBlank        = { E0},
    LcIdPersonalized = { F0}
  } lc_id_state_e;

  typedef enum logic [LcCountWidth-1:0] {
    LcCnt0  = {ZRO, ZRO, ZRO, ZRO, ZRO, ZRO, ZRO, ZRO, ZRO, ZRO, ZRO, ZRO, ZRO, ZRO, ZRO, ZRO},
    LcCnt1  = {C15, C14, C13, C12, C11, C10,  C9,  C8,  C7,  C6,  C5,  C4,  C3,  C2,  C1,  D0},
    LcCnt2  = {C15, C14, C13, C12, C11, C10,  C9,  C8,  C7,  C6,  C5,  C4,  C3,  C2,  D1,  D0},
    LcCnt3  = {C15, C14, C13, C12, C11, C10,  C9,  C8,  C7,  C6,  C5,  C4,  C3,  D2,  D1,  D0},
    LcCnt4  = {C15, C14, C13, C12, C11, C10,  C9,  C8,  C7,  C6,  C5,  C4,  D3,  D2,  D1,  D0},
    LcCnt5  = {C15, C14, C13, C12, C11, C10,  C9,  C8,  C7,  C6,  C5,  D4,  D3,  D2,  D1,  D0},
    LcCnt6  = {C15, C14, C13, C12, C11, C10,  C9,  C8,  C7,  C6,  D5,  D4,  D3,  D2,  D1,  D0},
    LcCnt7  = {C15, C14, C13, C12, C11, C10,  C9,  C8,  C7,  D6,  D5,  D4,  D3,  D2,  D1,  D0},
    LcCnt8  = {C15, C14, C13, C12, C11, C10,  C9,  C8,  D7,  D6,  D5,  D4,  D3,  D2,  D1,  D0},
    LcCnt9  = {C15, C14, C13, C12, C11, C10,  C9,  D8,  D7,  D6,  D5,  D4,  D3,  D2,  D1,  D0},
    LcCnt10 = {C15, C14, C13, C12, C11, C10,  D9,  D8,  D7,  D6,  D5,  D4,  D3,  D2,  D1,  D0},
    LcCnt11 = {C15, C14, C13, C12, C11, D10,  D9,  D8,  D7,  D6,  D5,  D4,  D3,  D2,  D1,  D0},
    LcCnt12 = {C15, C14, C13, C12, D11, D10,  D9,  D8,  D7,  D6,  D5,  D4,  D3,  D2,  D1,  D0},
    LcCnt13 = {C15, C14, C13, D12, D11, D10,  D9,  D8,  D7,  D6,  D5,  D4,  D3,  D2,  D1,  D0},
    LcCnt14 = {C15, C14, D13, D12, D11, D10,  D9,  D8,  D7,  D6,  D5,  D4,  D3,  D2,  D1,  D0},
    LcCnt15 = {C15, D14, D13, D12, D11, D10,  D9,  D8,  D7,  D6,  D5,  D4,  D3,  D2,  D1,  D0},
    LcCnt16 = {D15, D14, D13, D12, D11, D10,  D9,  D8,  D7,  D6,  D5,  D4,  D3,  D2,  D1,  D0}
  } lc_cnt_e;

  // Decoded life cycle state, used to interface with CSRs and TAP.
  typedef enum logic [DecLcStateWidth-1:0] {
    DecLcStRaw,
    DecLcStTestUnlocked0,
    DecLcStTestLocked0,
    DecLcStTestUnlocked1,
    DecLcStTestLocked1,
    DecLcStTestUnlocked2,
    DecLcStTestLocked2,
    DecLcStTestUnlocked3,
    DecLcStDev,
    DecLcStProd,
    DecLcStProdEnd,
    DecLcStRma,
    DecLcStScrap,
    DecLcStPostTrans,
    DecLcStEscalate,
    DecLcStInvalid
  } dec_lc_state_e;

  typedef enum logic [DecLcIdStateWidth-1:0] {
    DecLcIdBlank,
    DecLcIdPersonalized,
    DecLcIdInvalid
  } dec_lc_id_state_e;

  typedef logic [DecLcCountWidth-1:0] dec_lc_cnt_t;


  ///////////////////////////////////////////
  // Hashed RAW unlock and all-zero tokens //
  ///////////////////////////////////////////

  parameter int LcTokenWidth = 128;
  typedef logic [LcTokenWidth-1:0] lc_token_t;

  parameter lc_token_t AllZeroToken = {
    128'h0
  };
  parameter lc_token_t RndCnstRawUnlockToken = {
    128'h1C8BE2FF12790AE2E6D6A68151CBD084
  };
  parameter lc_token_t AllZeroTokenHashed = {
    128'h0
  };
  parameter lc_token_t RndCnstRawUnlockTokenHashed = {
    128'h1C8BE2FF12790AE2E6D6A68151CBD084
  };

endpackage : lc_ctrl_state_pkg


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//

package prim_ram_1p_pkg;

  typedef struct packed {
    logic       cfg_en;
    logic [3:0] cfg;
  } cfg_t;

  typedef struct packed {
    cfg_t ram_cfg;  // configuration for ram
    cfg_t rf_cfg;   // configuration for regfile
  } ram_1p_cfg_t;

  parameter ram_1p_cfg_t RAM_1P_CFG_DEFAULT = '0;

endpackage // prim_ram_1p_pkg

// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//

package lc_ctrl_pkg;

  import prim_util_pkg::vbits;
  import lc_ctrl_state_pkg::*;

  ///////////////////////////////////////
  // Netlist Constants (Hashed Tokens) //
  ///////////////////////////////////////

  parameter int NumTokens = 6;
  parameter int TokenIdxWidth = vbits(NumTokens);
  typedef enum logic [TokenIdxWidth-1:0] {
    // This is the index for the hashed all-zero constant.
    // All unconditional transitions use this token.
    ZeroTokenIdx       = 3'h0,
    RawUnlockTokenIdx  = 3'h1,
    TestUnlockTokenIdx = 3'h2,
    TestExitTokenIdx   = 3'h3,
    RmaTokenIdx        = 3'h4,
    // This is the index for an all-zero value (i.e., hashed value = '0).
    // This is used as an additional blocker for some invalid state transition edges.
    InvalidTokenIdx    = 3'h5
  } token_idx_e;

  ////////////////////////////////
  // Typedefs for LC Interfaces //
  ////////////////////////////////

  parameter int TxWidth = 4;

  typedef enum logic [TxWidth-1:0] {
    On  = 4'b1010,
    Off = 4'b0101
  } lc_tx_e;
  typedef logic [TxWidth-1:0] lc_tx_t;
  parameter lc_tx_t LC_TX_DEFAULT = lc_tx_t'(Off);

  parameter int RmaSeedWidth = 32;
  typedef logic [RmaSeedWidth-1:0] lc_flash_rma_seed_t;

  parameter int LcKeymgrDivWidth = 128;
  typedef logic [LcKeymgrDivWidth-1:0] lc_keymgr_div_t;

  ////////////////////
  // Main FSM State //
  ////////////////////

  // Encoding generated with:
  // $ ./sparse-fsm-encode.py -d 5 -m 14 -n 16 \
  //      -s 2934212379 --language=sv
  //
  // Hamming distance histogram:
  //
  //  0: --
  //  1: --
  //  2: --
  //  3: --
  //  4: --
  //  5: |||||| (6.59%)
  //  6: |||||||||| (10.99%)
  //  7: |||||||||||||||| (17.58%)
  //  8: |||||||||||||||||||| (20.88%)
  //  9: |||||||||||||||| (17.58%)
  // 10: |||||||||||||| (15.38%)
  // 11: |||||| (6.59%)
  // 12: ||| (3.30%)
  // 13: | (1.10%)
  // 14: --
  // 15: --
  // 16: --
  //
  // Minimum Hamming distance: 5
  // Maximum Hamming distance: 13
  //
  localparam int FsmStateWidth = 16;
  typedef enum logic [FsmStateWidth-1:0] {
    ResetSt       = 16'b1100000001111011,
    IdleSt        = 16'b1111011010111100,
    ClkMuxSt      = 16'b0000011110101101,
    CntIncrSt     = 16'b1100111011001001,
    CntProgSt     = 16'b0011001111000111,
    TransCheckSt  = 16'b0000110001010100,
    TokenHashSt   = 16'b1110100010001111,
    FlashRmaSt    = 16'b0110111010110000,
    TokenCheck0St = 16'b0010000011000000,
    TokenCheck1St = 16'b1101010101101111,
    TransProgSt   = 16'b1000000110101011,
    PostTransSt   = 16'b0110110100101100,
    EscalateSt    = 16'b1010100001010001,
    InvalidSt     = 16'b1011110110011011
  } fsm_state_e;

  ///////////////////////////////////////////
  // Manufacturing State Transition Matrix //
  ///////////////////////////////////////////

  // The token index matrix below encodes 1) which transition edges are valid and 2) which token
  // to use for a given transition edge. Note that unconditional but otherwise valid transitions
  // are assigned the ZeroTokenIdx, whereas invalid transitions are assigned an InvalidTokenIdx.
  parameter token_idx_e [NumLcStates-1:0][NumLcStates-1:0] TransTokenIdxMatrix = {
    // SCRAP
    {13{InvalidTokenIdx}}, // -> TEST_LOCKED0-2, TEST_UNLOCKED0-3, DEV, PROD, PROD_END, RMA, SCRAP
    // RMA
    ZeroTokenIdx,          // -> SCRAP
    {12{InvalidTokenIdx}}, // -> TEST_LOCKED0-2, TEST_UNLOCKED0-3, DEV, PROD, PROD_END, RMA
    // PROD_END
    ZeroTokenIdx,          // -> SCRAP
    {12{InvalidTokenIdx}}, // -> TEST_LOCKED0-2, TEST_UNLOCKED0-3, DEV, PROD, PROD_END, RMA
    // PROD
    ZeroTokenIdx,          // -> SCRAP
    RmaTokenIdx,           // -> RMA
    {11{InvalidTokenIdx}}, // -> TEST_LOCKED0-2, TEST_UNLOCKED0-3, DEV, PROD, PROD_END
    // DEV
    ZeroTokenIdx,          // -> SCRAP
    RmaTokenIdx,           // -> RMA
    {11{InvalidTokenIdx}}, // -> TEST_LOCKED0-2, TEST_UNLOCKED0-3, DEV, PROD, PROD_END
    // TEST_UNLOCKED3
    {2{ZeroTokenIdx}},     // -> SCRAP, RMA
    {3{TestExitTokenIdx}}, // -> PROD, PROD_END, DEV
    {8{InvalidTokenIdx}},  // -> TEST_LOCKED0-2, TEST_UNLOCKED0-3, RAW
    // TEST_LOCKED2
    ZeroTokenIdx,          // -> SCRAP
    InvalidTokenIdx,       // -> RMA
    {3{TestExitTokenIdx}}, // -> PROD, PROD_END, DEV
    TestUnlockTokenIdx,    // -> TEST_UNLOCKED3
    {7{InvalidTokenIdx}},  // -> TEST_LOCKED0-2, TEST_UNLOCKED0-2, RAW
    // TEST_UNLOCKED2
    {2{ZeroTokenIdx}},     // -> SCRAP, RMA
    {3{TestExitTokenIdx}}, // -> PROD, PROD_END, DEV
    InvalidTokenIdx,       // -> TEST_UNLOCKED3
    ZeroTokenIdx,          // -> TEST_LOCKED2
    {6{InvalidTokenIdx}},  // -> TEST_LOCKED0-1, TEST_UNLOCKED0-2, RAW
    // TEST_LOCKED1
    ZeroTokenIdx,          // -> SCRAP
    InvalidTokenIdx,       // -> RMA
    {3{TestExitTokenIdx}}, // -> PROD, PROD_END, DEV
    TestUnlockTokenIdx,    // -> TEST_UNLOCKED3
    InvalidTokenIdx  ,     // -> TEST_LOCKED2
    TestUnlockTokenIdx,    // -> TEST_UNLOCKED2
    {5{InvalidTokenIdx}},  // -> TEST_LOCKED0-1, TEST_UNLOCKED0-1, RAW
    // TEST_UNLOCKED1
    {2{ZeroTokenIdx}},     // -> SCRAP, RMA
    {3{TestExitTokenIdx}}, // -> PROD, PROD_END, DEV
    InvalidTokenIdx,       // -> TEST_UNLOCKED3
    ZeroTokenIdx,          // -> TEST_LOCKED2
    InvalidTokenIdx,       // -> TEST_UNLOCKED2
    ZeroTokenIdx,          // -> TEST_LOCKED1
    {4{InvalidTokenIdx}},  // -> TEST_LOCKED0, TEST_UNLOCKED0-1, RAW
    // TEST_LOCKED0
    ZeroTokenIdx,          // -> SCRAP
    InvalidTokenIdx,       // -> RMA
    {3{TestExitTokenIdx}}, // -> PROD, PROD_END, DEV
    TestUnlockTokenIdx,    // -> TEST_UNLOCKED3
    InvalidTokenIdx,       // -> TEST_LOCKED2
    TestUnlockTokenIdx,    // -> TEST_UNLOCKED2
    InvalidTokenIdx,       // -> TEST_LOCKED1
    TestUnlockTokenIdx,    // -> TEST_UNLOCKED1
    {3{InvalidTokenIdx}},  // -> TEST_LOCKED0, TEST_UNLOCKED0, RAW
    // TEST_UNLOCKED0
    {2{ZeroTokenIdx}},     // -> SCRAP, RMA
    {3{TestExitTokenIdx}}, // -> PROD, PROD_END, DEV
    InvalidTokenIdx,       // -> TEST_UNLOCKED3
    ZeroTokenIdx,          // -> TEST_LOCKED2
    InvalidTokenIdx,       // -> TEST_UNLOCKED2
    ZeroTokenIdx,          // -> TEST_LOCKED1
    InvalidTokenIdx,       // -> TEST_UNLOCKED1
    ZeroTokenIdx,          // -> TEST_LOCKED0
    {2{InvalidTokenIdx}},  // -> TEST_UNLOCKED0, RAW
    // RAW
    ZeroTokenIdx,          // -> SCRAP
    {4{InvalidTokenIdx}},  // -> RMA, PROD, PROD_END, DEV
    RawUnlockTokenIdx,     // -> TEST_UNLOCKED3
    InvalidTokenIdx,       // -> TEST_LOCKED2
    RawUnlockTokenIdx,     // -> TEST_UNLOCKED2
    InvalidTokenIdx,       // -> TEST_LOCKED1
    RawUnlockTokenIdx,     // -> TEST_UNLOCKED1
    InvalidTokenIdx,       // -> TEST_LOCKED0
    RawUnlockTokenIdx,     // -> TEST_UNLOCKED0
    InvalidTokenIdx        // -> RAW
  };

endpackage : lc_ctrl_pkg

// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

package prim_esc_pkg;

  typedef struct packed {
    logic esc_p;
    logic esc_n;
  } esc_tx_t;

  typedef struct packed {
    logic resp_p;
    logic resp_n;
  } esc_rx_t;

  parameter esc_tx_t ESC_TX_DEFAULT = '{esc_p:  1'b0,
                                        esc_n:  1'b1};

  parameter esc_rx_t ESC_RX_DEFAULT = '{resp_p: 1'b0,
                                        resp_n: 1'b1};

endpackage : prim_esc_pkg


module paramod00798253a2da2b158adcde19e501253b4257bf48auxy_ibex_core (clk_i, rst_ni, hart_id_i, boot_addr_i, instr_req_o, instr_gnt_i, instr_rvalid_i, instr_addr_o, instr_rdata_i, instr_err_i, data_req_o, data_gnt_i, data_rvalid_i, data_we_o, data_be_o, data_addr_o, data_wdata_o, data_rdata_i, data_err_i, dummy_instr_id_o, rf_raddr_a_o
, rf_raddr_b_o, rf_waddr_wb_o, rf_we_wb_o, rf_wdata_wb_ecc_o, rf_rdata_a_ecc_i, rf_rdata_b_ecc_i, ic_tag_req_o, ic_tag_write_o, ic_tag_addr_o, ic_tag_wdata_o, ic_tag_rdata_i, ic_data_req_o, ic_data_write_o, ic_data_addr_o, ic_data_wdata_o, ic_data_rdata_i, irq_software_i, irq_timer_i, irq_external_i, irq_fast_i, irq_nm_i
, irq_pending_o, debug_req_i, crash_dump_o, alert_minor_o, alert_major_o, core_busy_o, ic_tag_write_o_t0, ic_tag_wdata_o_t0, ic_tag_req_o_t0, ic_tag_rdata_i_t0, ic_tag_addr_o_t0, ic_data_write_o_t0, ic_data_wdata_o_t0, ic_data_req_o_t0, ic_data_rdata_i_t0, ic_data_addr_o_t0, boot_addr_i_t0, dummy_instr_id_o_t0, instr_rvalid_i_t0, instr_req_o_t0, instr_rdata_i_t0
, instr_gnt_i_t0, instr_err_i_t0, instr_addr_o_t0, data_req_o_t0, rf_raddr_a_o_t0, rf_raddr_b_o_t0, data_we_o_t0, debug_req_i_t0, irq_nm_i_t0, data_addr_o_t0, data_be_o_t0, data_err_i_t0, data_gnt_i_t0, data_rdata_i_t0, data_rvalid_i_t0, data_wdata_o_t0, rf_waddr_wb_o_t0, rf_we_wb_o_t0, hart_id_i_t0, irq_external_i_t0, irq_fast_i_t0
, irq_pending_o_t0, irq_software_i_t0, irq_timer_i_t0, alert_major_o_t0, alert_minor_o_t0, core_busy_o_t0, crash_dump_o_t0, rf_rdata_a_ecc_i_t0, rf_rdata_b_ecc_i_t0, rf_wdata_wb_ecc_o_t0);
  wire _00_;
  wire _01_;
  wire _02_;
  wire _03_;
  wire _04_;
  wire _05_;
  wire _06_;
  wire _07_;
  wire [11:0] _08_;
  wire _09_;
  wire _10_;
  wire _11_;
  wire _12_;
  wire _13_;
  wire _14_;
  wire _15_;
  wire _16_;
  wire _17_;
  wire _18_;
  wire _19_;
  wire _20_;
  wire _21_;
  wire _22_;
  wire _23_;
  wire [11:0] _24_;
  wire [11:0] _25_;
  wire [11:0] _26_;
  wire _27_;
  wire _28_;
  wire _29_;
  wire _30_;
  wire _31_;
  wire [11:0] _32_;
  wire [11:0] _33_;
  wire [11:0] _34_;
  wire _35_;
  wire _36_;
  wire _37_;
  output alert_major_o;
  wire alert_major_o;
  output alert_major_o_t0;
  wire alert_major_o_t0;
  output alert_minor_o;
  wire alert_minor_o;
  output alert_minor_o_t0;
  wire alert_minor_o_t0;
  wire [31:0] alu_adder_result_ex;
  wire [31:0] alu_adder_result_ex_t0;
  wire [31:0] alu_operand_a_ex;
  wire [31:0] alu_operand_a_ex_t0;
  wire [31:0] alu_operand_b_ex;
  wire [31:0] alu_operand_b_ex_t0;
  wire [5:0] alu_operator_ex;
  wire [5:0] alu_operator_ex_t0;
  input [31:0] boot_addr_i;
  wire [31:0] boot_addr_i;
  input [31:0] boot_addr_i_t0;
  wire [31:0] boot_addr_i_t0;
  wire branch_decision;
  wire branch_decision_t0;
  wire [31:0] branch_target_ex;
  wire [31:0] branch_target_ex_t0;
  wire [31:0] bt_a_operand;
  wire [31:0] bt_a_operand_t0;
  wire [31:0] bt_b_operand;
  wire [31:0] bt_b_operand_t0;
  input clk_i;
  wire clk_i;
  output core_busy_o;
  wire core_busy_o;
  output core_busy_o_t0;
  wire core_busy_o_t0;
  output [127:0] crash_dump_o;
  wire [127:0] crash_dump_o;
  output [127:0] crash_dump_o_t0;
  wire [127:0] crash_dump_o_t0;
  wire csr_access;
  wire csr_access_t0;
  wire [11:0] csr_addr;
  wire [11:0] csr_addr_t0;
  wire [31:0] csr_depc;
  wire [31:0] csr_depc_t0;
  wire [31:0] csr_mepc;
  wire [31:0] csr_mepc_t0;
  wire csr_mstatus_mie;
  wire csr_mstatus_mie_t0;
  wire csr_mstatus_tw;
  wire csr_mstatus_tw_t0;
  wire [31:0] csr_mtval;
  wire [31:0] csr_mtval_t0;
  wire [31:0] csr_mtvec;
  wire csr_mtvec_init;
  wire csr_mtvec_init_t0;
  wire [31:0] csr_mtvec_t0;
  wire [1:0] csr_op;
  wire csr_op_en;
  wire csr_op_en_t0;
  wire [1:0] csr_op_t0;
  wire [135:0] csr_pmp_addr;
  wire [135:0] csr_pmp_addr_t0;
  wire [23:0] csr_pmp_cfg;
  wire [23:0] csr_pmp_cfg_t0;
  wire [2:0] csr_pmp_mseccfg;
  wire [2:0] csr_pmp_mseccfg_t0;
  wire [31:0] csr_rdata;
  wire [31:0] csr_rdata_t0;
  wire csr_restore_dret_id;
  wire csr_restore_dret_id_t0;
  wire csr_restore_mret_id;
  wire csr_restore_mret_id_t0;
  wire csr_save_cause;
  wire csr_save_cause_t0;
  wire csr_save_id;
  wire csr_save_id_t0;
  wire csr_save_if;
  wire csr_save_if_t0;
  wire csr_save_wb;
  wire csr_save_wb_t0;
  wire csr_shadow_err;
  wire csr_shadow_err_t0;
  wire ctrl_busy;
  wire ctrl_busy_t0;
  output [31:0] data_addr_o;
  wire [31:0] data_addr_o;
  output [31:0] data_addr_o_t0;
  wire [31:0] data_addr_o_t0;
  output [3:0] data_be_o;
  wire [3:0] data_be_o;
  output [3:0] data_be_o_t0;
  wire [3:0] data_be_o_t0;
  input data_err_i;
  wire data_err_i;
  input data_err_i_t0;
  wire data_err_i_t0;
  input data_gnt_i;
  wire data_gnt_i;
  input data_gnt_i_t0;
  wire data_gnt_i_t0;
  wire data_ind_timing;
  wire data_ind_timing_t0;
  input [31:0] data_rdata_i;
  wire [31:0] data_rdata_i;
  input [31:0] data_rdata_i_t0;
  wire [31:0] data_rdata_i_t0;
  output data_req_o;
  wire data_req_o;
  output data_req_o_t0;
  wire data_req_o_t0;
  input data_rvalid_i;
  wire data_rvalid_i;
  input data_rvalid_i_t0;
  wire data_rvalid_i_t0;
  output [31:0] data_wdata_o;
  wire [31:0] data_wdata_o;
  output [31:0] data_wdata_o_t0;
  wire [31:0] data_wdata_o_t0;
  output data_we_o;
  wire data_we_o;
  output data_we_o_t0;
  wire data_we_o_t0;
  wire [2:0] debug_cause;
  wire [2:0] debug_cause_t0;
  wire debug_csr_save;
  wire debug_csr_save_t0;
  wire debug_ebreakm;
  wire debug_ebreakm_t0;
  wire debug_ebreaku;
  wire debug_ebreaku_t0;
  wire debug_mode;
  wire debug_mode_t0;
  input debug_req_i;
  wire debug_req_i;
  input debug_req_i_t0;
  wire debug_req_i_t0;
  wire debug_single_step;
  wire debug_single_step_t0;
  wire div_en_ex;
  wire div_en_ex_t0;
  wire div_sel_ex;
  wire div_sel_ex_t0;
  wire dummy_instr_en;
  wire dummy_instr_en_t0;
  output dummy_instr_id_o;
  wire dummy_instr_id_o;
  output dummy_instr_id_o_t0;
  wire dummy_instr_id_o_t0;
  wire [2:0] dummy_instr_mask;
  wire [2:0] dummy_instr_mask_t0;
  wire [31:0] dummy_instr_seed;
  wire dummy_instr_seed_en;
  wire dummy_instr_seed_en_t0;
  wire [31:0] dummy_instr_seed_t0;
  wire en_wb;
  wire en_wb_t0;
  wire ex_valid;
  wire ex_valid_t0;
  wire [5:0] exc_cause;
  wire [5:0] exc_cause_t0;
  wire [1:0] exc_pc_mux_id;
  wire [1:0] exc_pc_mux_id_t0;
  wire [1:0] \g_no_pmp.unused_priv_lvl_if ;
  wire [1:0] \g_no_pmp.unused_priv_lvl_if_t0 ;
  wire [1:0] \g_no_pmp.unused_priv_lvl_ls ;
  wire [1:0] \g_no_pmp.unused_priv_lvl_ls_t0 ;
  wire \gen_no_regfile_ecc.unused_rf_rd_a_wb_match ;
  wire \gen_no_regfile_ecc.unused_rf_rd_a_wb_match_t0 ;
  wire \gen_no_regfile_ecc.unused_rf_rd_b_wb_match ;
  wire \gen_no_regfile_ecc.unused_rf_rd_b_wb_match_t0 ;
  wire \gen_no_regfile_ecc.unused_rf_ren_a ;
  wire \gen_no_regfile_ecc.unused_rf_ren_a_t0 ;
  wire \gen_no_regfile_ecc.unused_rf_ren_b ;
  wire \gen_no_regfile_ecc.unused_rf_ren_b_t0 ;
  input [31:0] hart_id_i;
  wire [31:0] hart_id_i;
  input [31:0] hart_id_i_t0;
  wire [31:0] hart_id_i_t0;
  output [7:0] ic_data_addr_o;
  wire [7:0] ic_data_addr_o;
  output [7:0] ic_data_addr_o_t0;
  wire [7:0] ic_data_addr_o_t0;
  input [127:0] ic_data_rdata_i;
  wire [127:0] ic_data_rdata_i;
  input [127:0] ic_data_rdata_i_t0;
  wire [127:0] ic_data_rdata_i_t0;
  output [1:0] ic_data_req_o;
  wire [1:0] ic_data_req_o;
  output [1:0] ic_data_req_o_t0;
  wire [1:0] ic_data_req_o_t0;
  output [63:0] ic_data_wdata_o;
  wire [63:0] ic_data_wdata_o;
  output [63:0] ic_data_wdata_o_t0;
  wire [63:0] ic_data_wdata_o_t0;
  output ic_data_write_o;
  wire ic_data_write_o;
  output ic_data_write_o_t0;
  wire ic_data_write_o_t0;
  output [7:0] ic_tag_addr_o;
  wire [7:0] ic_tag_addr_o;
  output [7:0] ic_tag_addr_o_t0;
  wire [7:0] ic_tag_addr_o_t0;
  input [43:0] ic_tag_rdata_i;
  wire [43:0] ic_tag_rdata_i;
  input [43:0] ic_tag_rdata_i_t0;
  wire [43:0] ic_tag_rdata_i_t0;
  output [1:0] ic_tag_req_o;
  wire [1:0] ic_tag_req_o;
  output [1:0] ic_tag_req_o_t0;
  wire [1:0] ic_tag_req_o_t0;
  output [21:0] ic_tag_wdata_o;
  wire [21:0] ic_tag_wdata_o;
  output [21:0] ic_tag_wdata_o_t0;
  wire [21:0] ic_tag_wdata_o_t0;
  output ic_tag_write_o;
  wire ic_tag_write_o;
  output ic_tag_write_o_t0;
  wire ic_tag_write_o_t0;
  wire icache_enable;
  wire icache_enable_t0;
  wire icache_inval;
  wire icache_inval_t0;
  wire id_in_ready;
  wire id_in_ready_t0;
  wire if_busy;
  wire if_busy_t0;
  wire illegal_c_insn_id;
  wire illegal_c_insn_id_t0;
  wire illegal_csr_insn_id;
  wire illegal_csr_insn_id_t0;
  wire illegal_insn_id;
  wire illegal_insn_id_t0;
  wire [67:0] imd_val_d_ex;
  wire [67:0] imd_val_d_ex_t0;
  wire [67:0] imd_val_q_ex;
  wire [67:0] imd_val_q_ex_t0;
  wire [1:0] imd_val_we_ex;
  wire [1:0] imd_val_we_ex_t0;
  output [31:0] instr_addr_o;
  wire [31:0] instr_addr_o;
  output [31:0] instr_addr_o_t0;
  wire [31:0] instr_addr_o_t0;
  wire instr_bp_taken_id;
  wire instr_bp_taken_id_t0;
  wire instr_done_wb;
  wire instr_done_wb_t0;
  input instr_err_i;
  wire instr_err_i;
  input instr_err_i_t0;
  wire instr_err_i_t0;
  wire instr_fetch_err;
  wire instr_fetch_err_plus2;
  wire instr_fetch_err_plus2_t0;
  wire instr_fetch_err_t0;
  wire instr_first_cycle_id;
  wire instr_first_cycle_id_t0;
  input instr_gnt_i;
  wire instr_gnt_i;
  input instr_gnt_i_t0;
  wire instr_gnt_i_t0;
  wire instr_id_done;
  wire instr_id_done_t0;
  wire instr_is_compressed_id;
  wire instr_is_compressed_id_t0;
  wire instr_new_id;
  wire instr_new_id_t0;
  wire instr_perf_count_id;
  wire instr_perf_count_id_t0;
  wire [31:0] instr_rdata_alu_id;
  wire [31:0] instr_rdata_alu_id_t0;
  wire [15:0] instr_rdata_c_id;
  wire [15:0] instr_rdata_c_id_t0;
  input [31:0] instr_rdata_i;
  wire [31:0] instr_rdata_i;
  input [31:0] instr_rdata_i_t0;
  wire [31:0] instr_rdata_i_t0;
  wire [31:0] instr_rdata_id;
  wire [31:0] instr_rdata_id_t0;
  wire instr_req_int;
  wire instr_req_int_t0;
  output instr_req_o;
  wire instr_req_o;
  output instr_req_o_t0;
  wire instr_req_o_t0;
  input instr_rvalid_i;
  wire instr_rvalid_i;
  input instr_rvalid_i_t0;
  wire instr_rvalid_i_t0;
  wire [1:0] instr_type_wb;
  wire [1:0] instr_type_wb_t0;
  wire instr_valid_clear;
  wire instr_valid_clear_t0;
  wire instr_valid_id;
  wire instr_valid_id_t0;
  input irq_external_i;
  wire irq_external_i;
  input irq_external_i_t0;
  wire irq_external_i_t0;
  input [14:0] irq_fast_i;
  wire [14:0] irq_fast_i;
  input [14:0] irq_fast_i_t0;
  wire [14:0] irq_fast_i_t0;
  input irq_nm_i;
  wire irq_nm_i;
  input irq_nm_i_t0;
  wire irq_nm_i_t0;
  output irq_pending_o;
  wire irq_pending_o;
  output irq_pending_o_t0;
  wire irq_pending_o_t0;
  input irq_software_i;
  wire irq_software_i;
  input irq_software_i_t0;
  wire irq_software_i_t0;
  input irq_timer_i;
  wire irq_timer_i;
  input irq_timer_i_t0;
  wire irq_timer_i_t0;
  wire [17:0] irqs;
  wire [17:0] irqs_t0;
  wire lsu_addr_incr_req;
  wire lsu_addr_incr_req_t0;
  wire [31:0] lsu_addr_last;
  wire [31:0] lsu_addr_last_t0;
  wire lsu_busy;
  wire lsu_busy_t0;
  wire lsu_load_err;
  wire lsu_load_err_t0;
  wire lsu_req;
  wire lsu_req_done;
  wire lsu_req_done_t0;
  wire lsu_req_t0;
  wire lsu_resp_err;
  wire lsu_resp_err_t0;
  wire lsu_resp_valid;
  wire lsu_resp_valid_t0;
  wire lsu_sign_ext;
  wire lsu_sign_ext_t0;
  wire lsu_store_err;
  wire lsu_store_err_t0;
  wire [1:0] lsu_type;
  wire [1:0] lsu_type_t0;
  wire [31:0] lsu_wdata;
  wire [31:0] lsu_wdata_t0;
  wire lsu_we;
  wire lsu_we_t0;
  wire mult_en_ex;
  wire mult_en_ex_t0;
  wire mult_sel_ex;
  wire mult_sel_ex_t0;
  wire [31:0] multdiv_operand_a_ex;
  wire [31:0] multdiv_operand_a_ex_t0;
  wire [31:0] multdiv_operand_b_ex;
  wire [31:0] multdiv_operand_b_ex_t0;
  wire [1:0] multdiv_operator_ex;
  wire [1:0] multdiv_operator_ex_t0;
  wire multdiv_ready_id;
  wire multdiv_ready_id_t0;
  wire [1:0] multdiv_signed_mode_ex;
  wire [1:0] multdiv_signed_mode_ex_t0;
  wire nmi_mode;
  wire nmi_mode_t0;
  wire nt_branch_mispredict;
  wire nt_branch_mispredict_t0;
  wire outstanding_load_wb;
  wire outstanding_load_wb_t0;
  wire outstanding_store_wb;
  wire outstanding_store_wb_t0;
  wire [31:0] pc_id /* verilator public */;
  wire [31:0] pc_id_t0 /* verilator public */;
  wire [31:0] pc_if;
  wire [31:0] pc_if_t0;
  wire pc_mismatch_alert;
  wire pc_mismatch_alert_t0;
  wire [2:0] pc_mux_id;
  wire [2:0] pc_mux_id_t0;
  wire pc_set;
  wire pc_set_spec;
  wire pc_set_spec_t0;
  wire pc_set_t0;
  wire [31:0] pc_wb;
  wire [31:0] pc_wb_t0;
  wire perf_branch;
  wire perf_branch_t0;
  wire perf_div_wait;
  wire perf_div_wait_t0;
  wire perf_dside_wait;
  wire perf_dside_wait_t0;
  wire perf_instr_ret_compressed_wb;
  wire perf_instr_ret_compressed_wb_t0;
  wire perf_instr_ret_wb;
  wire perf_instr_ret_wb_t0;
  wire perf_iside_wait;
  wire perf_iside_wait_t0;
  wire perf_jump;
  wire perf_jump_t0;
  wire perf_load;
  wire perf_load_t0;
  wire perf_mul_wait;
  wire perf_mul_wait_t0;
  wire perf_store;
  wire perf_store_t0;
  wire perf_tbranch;
  wire perf_tbranch_t0;
  wire [1:0] priv_mode_id;
  wire [1:0] priv_mode_id_t0;
  wire ready_wb;
  wire ready_wb_t0;
  wire [31:0] result_ex;
  wire [31:0] result_ex_t0;
  output [4:0] rf_raddr_a_o;
  wire [4:0] rf_raddr_a_o;
  output [4:0] rf_raddr_a_o_t0;
  wire [4:0] rf_raddr_a_o_t0;
  output [4:0] rf_raddr_b_o;
  wire [4:0] rf_raddr_b_o;
  output [4:0] rf_raddr_b_o_t0;
  wire [4:0] rf_raddr_b_o_t0;
  input [31:0] rf_rdata_a_ecc_i;
  wire [31:0] rf_rdata_a_ecc_i;
  input [31:0] rf_rdata_a_ecc_i_t0;
  wire [31:0] rf_rdata_a_ecc_i_t0;
  input [31:0] rf_rdata_b_ecc_i;
  wire [31:0] rf_rdata_b_ecc_i;
  input [31:0] rf_rdata_b_ecc_i_t0;
  wire [31:0] rf_rdata_b_ecc_i_t0;
  wire [4:0] rf_waddr_id;
  wire [4:0] rf_waddr_id_t0;
  output [4:0] rf_waddr_wb_o;
  wire [4:0] rf_waddr_wb_o;
  output [4:0] rf_waddr_wb_o_t0;
  wire [4:0] rf_waddr_wb_o_t0;
  wire [31:0] rf_wdata_fwd_wb;
  wire [31:0] rf_wdata_fwd_wb_t0;
  wire [31:0] rf_wdata_id;
  wire [31:0] rf_wdata_id_t0;
  wire [31:0] rf_wdata_lsu;
  wire [31:0] rf_wdata_lsu_t0;
  output [31:0] rf_wdata_wb_ecc_o;
  wire [31:0] rf_wdata_wb_ecc_o;
  output [31:0] rf_wdata_wb_ecc_o_t0;
  wire [31:0] rf_wdata_wb_ecc_o_t0;
  wire rf_we_id;
  wire rf_we_id_t0;
  wire rf_we_lsu;
  wire rf_we_lsu_t0;
  output rf_we_wb_o;
  wire rf_we_wb_o;
  output rf_we_wb_o_t0;
  wire rf_we_wb_o_t0;
  wire rf_write_wb;
  wire rf_write_wb_t0;
  input rst_ni;
  wire rst_ni;
  wire trigger_match;
  wire trigger_match_t0;
  assign perf_iside_wait = id_in_ready & _35_;
  assign _09_ = id_in_ready_t0 & _35_;
  assign _10_ = instr_valid_id_t0 & id_in_ready;
  assign _11_ = id_in_ready_t0 & instr_valid_id_t0;
  assign _27_ = _09_ | _10_;
  assign perf_iside_wait_t0 = _27_ | _11_;
  assign _08_ = ~ { csr_access, csr_access, csr_access, csr_access, csr_access, csr_access, csr_access, csr_access, csr_access, csr_access, csr_access, csr_access };
  assign _32_ = { csr_access_t0, csr_access_t0, csr_access_t0, csr_access_t0, csr_access_t0, csr_access_t0, csr_access_t0, csr_access_t0, csr_access_t0, csr_access_t0, csr_access_t0, csr_access_t0 } | _08_;
  assign _33_ = { csr_access_t0, csr_access_t0, csr_access_t0, csr_access_t0, csr_access_t0, csr_access_t0, csr_access_t0, csr_access_t0, csr_access_t0, csr_access_t0, csr_access_t0, csr_access_t0 } | { csr_access, csr_access, csr_access, csr_access, csr_access, csr_access, csr_access, csr_access, csr_access, csr_access, csr_access, csr_access };
  assign _24_ = 12'h000 & _32_;
  assign _25_ = alu_operand_b_ex_t0[11:0] & _33_;
  assign _34_ = _24_ | _25_;
  assign _26_ = { csr_access_t0, csr_access_t0, csr_access_t0, csr_access_t0, csr_access_t0, csr_access_t0, csr_access_t0, csr_access_t0, csr_access_t0, csr_access_t0, csr_access_t0, csr_access_t0 } & alu_operand_b_ex[11:0];
  assign csr_addr_t0 = _26_ | _34_;
  assign _00_ = ~ ctrl_busy;
  assign _02_ = ~ _36_;
  assign _04_ = ~ lsu_load_err;
  assign _06_ = ~ pc_mismatch_alert;
  assign _01_ = ~ if_busy;
  assign _03_ = ~ lsu_busy;
  assign _05_ = ~ lsu_store_err;
  assign _07_ = ~ csr_shadow_err;
  assign _12_ = ctrl_busy_t0 & _01_;
  assign _15_ = _37_ & _03_;
  assign _18_ = lsu_load_err_t0 & _05_;
  assign _21_ = pc_mismatch_alert_t0 & _07_;
  assign _13_ = if_busy_t0 & _00_;
  assign _16_ = lsu_busy_t0 & _02_;
  assign _19_ = lsu_store_err_t0 & _04_;
  assign _22_ = csr_shadow_err_t0 & _06_;
  assign _14_ = ctrl_busy_t0 & if_busy_t0;
  assign _17_ = _37_ & lsu_busy_t0;
  assign _20_ = lsu_load_err_t0 & lsu_store_err_t0;
  assign _23_ = pc_mismatch_alert_t0 & csr_shadow_err_t0;
  assign _28_ = _12_ | _13_;
  assign _29_ = _15_ | _16_;
  assign _30_ = _18_ | _19_;
  assign _31_ = _21_ | _22_;
  assign _37_ = _28_ | _14_;
  assign core_busy_o_t0 = _29_ | _17_;
  assign lsu_resp_err_t0 = _30_ | _20_;
  assign alert_major_o_t0 = _31_ | _23_;
  assign _35_ = ~ instr_valid_id;
  assign _36_ = ctrl_busy | if_busy;
  assign core_busy_o = _36_ | lsu_busy;
  assign lsu_resp_err = lsu_load_err | lsu_store_err;
  assign alert_major_o = pc_mismatch_alert | csr_shadow_err;
  assign csr_addr = csr_access ? alu_operand_b_ex[11:0] : 12'h000;
  paramoda7b3f37e1f713a4d0901b62b3f601f61ae6218e0auxy_ibex_cs_registers  cs_registers_i (
    .boot_addr_i(boot_addr_i),
    .boot_addr_i_t0(boot_addr_i_t0),
    .branch_i(perf_branch),
    .branch_i_t0(perf_branch_t0),
    .branch_taken_i(perf_tbranch),
    .branch_taken_i_t0(perf_tbranch_t0),
    .clk_i(clk_i),
    .csr_access_i(csr_access),
    .csr_access_i_t0(csr_access_t0),
    .csr_addr_i(csr_addr),
    .csr_addr_i_t0(csr_addr_t0),
    .csr_depc_o(csr_depc),
    .csr_depc_o_t0(csr_depc_t0),
    .csr_mcause_i(exc_cause),
    .csr_mcause_i_t0(exc_cause_t0),
    .csr_mepc_o(csr_mepc),
    .csr_mepc_o_t0(csr_mepc_t0),
    .csr_mstatus_mie_o(csr_mstatus_mie),
    .csr_mstatus_mie_o_t0(csr_mstatus_mie_t0),
    .csr_mstatus_tw_o(csr_mstatus_tw),
    .csr_mstatus_tw_o_t0(csr_mstatus_tw_t0),
    .csr_mtval_i(csr_mtval),
    .csr_mtval_i_t0(csr_mtval_t0),
    .csr_mtvec_init_i(csr_mtvec_init),
    .csr_mtvec_init_i_t0(csr_mtvec_init_t0),
    .csr_mtvec_o(csr_mtvec),
    .csr_mtvec_o_t0(csr_mtvec_t0),
    .csr_op_en_i(csr_op_en),
    .csr_op_en_i_t0(csr_op_en_t0),
    .csr_op_i(csr_op),
    .csr_op_i_t0(csr_op_t0),
    .csr_pmp_addr_o(csr_pmp_addr),
    .csr_pmp_addr_o_t0(csr_pmp_addr_t0),
    .csr_pmp_cfg_o(csr_pmp_cfg),
    .csr_pmp_cfg_o_t0(csr_pmp_cfg_t0),
    .csr_pmp_mseccfg_o(csr_pmp_mseccfg),
    .csr_pmp_mseccfg_o_t0(csr_pmp_mseccfg_t0),
    .csr_rdata_o(csr_rdata),
    .csr_rdata_o_t0(csr_rdata_t0),
    .csr_restore_dret_i(csr_restore_dret_id),
    .csr_restore_dret_i_t0(csr_restore_dret_id_t0),
    .csr_restore_mret_i(csr_restore_mret_id),
    .csr_restore_mret_i_t0(csr_restore_mret_id_t0),
    .csr_save_cause_i(csr_save_cause),
    .csr_save_cause_i_t0(csr_save_cause_t0),
    .csr_save_id_i(csr_save_id),
    .csr_save_id_i_t0(csr_save_id_t0),
    .csr_save_if_i(csr_save_if),
    .csr_save_if_i_t0(csr_save_if_t0),
    .csr_save_wb_i(csr_save_wb),
    .csr_save_wb_i_t0(csr_save_wb_t0),
    .csr_shadow_err_o(csr_shadow_err),
    .csr_shadow_err_o_t0(csr_shadow_err_t0),
    .csr_wdata_i(alu_operand_a_ex),
    .csr_wdata_i_t0(alu_operand_a_ex_t0),
    .data_ind_timing_o(data_ind_timing),
    .data_ind_timing_o_t0(data_ind_timing_t0),
    .debug_cause_i(debug_cause),
    .debug_cause_i_t0(debug_cause_t0),
    .debug_csr_save_i(debug_csr_save),
    .debug_csr_save_i_t0(debug_csr_save_t0),
    .debug_ebreakm_o(debug_ebreakm),
    .debug_ebreakm_o_t0(debug_ebreakm_t0),
    .debug_ebreaku_o(debug_ebreaku),
    .debug_ebreaku_o_t0(debug_ebreaku_t0),
    .debug_mode_i(debug_mode),
    .debug_mode_i_t0(debug_mode_t0),
    .debug_single_step_o(debug_single_step),
    .debug_single_step_o_t0(debug_single_step_t0),
    .div_wait_i(perf_div_wait),
    .div_wait_i_t0(perf_div_wait_t0),
    .dside_wait_i(perf_dside_wait),
    .dside_wait_i_t0(perf_dside_wait_t0),
    .dummy_instr_en_o(dummy_instr_en),
    .dummy_instr_en_o_t0(dummy_instr_en_t0),
    .dummy_instr_mask_o(dummy_instr_mask),
    .dummy_instr_mask_o_t0(dummy_instr_mask_t0),
    .dummy_instr_seed_en_o(dummy_instr_seed_en),
    .dummy_instr_seed_en_o_t0(dummy_instr_seed_en_t0),
    .dummy_instr_seed_o(dummy_instr_seed),
    .dummy_instr_seed_o_t0(dummy_instr_seed_t0),
    .hart_id_i(hart_id_i),
    .hart_id_i_t0(hart_id_i_t0),
    .icache_enable_o(icache_enable),
    .icache_enable_o_t0(icache_enable_t0),
    .illegal_csr_insn_o(illegal_csr_insn_id),
    .illegal_csr_insn_o_t0(illegal_csr_insn_id_t0),
    .instr_ret_compressed_i(perf_instr_ret_compressed_wb),
    .instr_ret_compressed_i_t0(perf_instr_ret_compressed_wb_t0),
    .instr_ret_i(perf_instr_ret_wb),
    .instr_ret_i_t0(perf_instr_ret_wb_t0),
    .irq_external_i(irq_external_i),
    .irq_external_i_t0(irq_external_i_t0),
    .irq_fast_i(irq_fast_i),
    .irq_fast_i_t0(irq_fast_i_t0),
    .irq_pending_o(irq_pending_o),
    .irq_pending_o_t0(irq_pending_o_t0),
    .irq_software_i(irq_software_i),
    .irq_software_i_t0(irq_software_i_t0),
    .irq_timer_i(irq_timer_i),
    .irq_timer_i_t0(irq_timer_i_t0),
    .irqs_o(irqs),
    .irqs_o_t0(irqs_t0),
    .iside_wait_i(perf_iside_wait),
    .iside_wait_i_t0(perf_iside_wait_t0),
    .jump_i(perf_jump),
    .jump_i_t0(perf_jump_t0),
    .mem_load_i(perf_load),
    .mem_load_i_t0(perf_load_t0),
    .mem_store_i(perf_store),
    .mem_store_i_t0(perf_store_t0),
    .mul_wait_i(perf_mul_wait),
    .mul_wait_i_t0(perf_mul_wait_t0),
    .nmi_mode_i(nmi_mode),
    .nmi_mode_i_t0(nmi_mode_t0),
    .pc_id_i(pc_id),
    .pc_id_i_t0(pc_id_t0),
    .pc_if_i(pc_if),
    .pc_if_i_t0(pc_if_t0),
    .pc_wb_i(pc_wb),
    .pc_wb_i_t0(pc_wb_t0),
    .priv_mode_id_o(priv_mode_id),
    .priv_mode_id_o_t0(priv_mode_id_t0),
    .priv_mode_if_o(\g_no_pmp.unused_priv_lvl_if ),
    .priv_mode_if_o_t0(\g_no_pmp.unused_priv_lvl_if_t0 ),
    .priv_mode_lsu_o(\g_no_pmp.unused_priv_lvl_ls ),
    .priv_mode_lsu_o_t0(\g_no_pmp.unused_priv_lvl_ls_t0 ),
    .rst_ni(rst_ni),
    .trigger_match_o(trigger_match),
    .trigger_match_o_t0(trigger_match_t0)
  );
  paramodc28f38d36bce0367a978a541cbb5da157ce66eceauxy_ibex_ex_block  ex_block_i (
    .alu_adder_result_ex_o(alu_adder_result_ex),
    .alu_adder_result_ex_o_t0(alu_adder_result_ex_t0),
    .alu_instr_first_cycle_i(instr_first_cycle_id),
    .alu_instr_first_cycle_i_t0(instr_first_cycle_id_t0),
    .alu_operand_a_i(alu_operand_a_ex),
    .alu_operand_a_i_t0(alu_operand_a_ex_t0),
    .alu_operand_b_i(alu_operand_b_ex),
    .alu_operand_b_i_t0(alu_operand_b_ex_t0),
    .alu_operator_i(alu_operator_ex),
    .alu_operator_i_t0(alu_operator_ex_t0),
    .branch_decision_o(branch_decision),
    .branch_decision_o_t0(branch_decision_t0),
    .branch_target_o(branch_target_ex),
    .branch_target_o_t0(branch_target_ex_t0),
    .bt_a_operand_i(bt_a_operand),
    .bt_a_operand_i_t0(bt_a_operand_t0),
    .bt_b_operand_i(bt_b_operand),
    .bt_b_operand_i_t0(bt_b_operand_t0),
    .clk_i(clk_i),
    .data_ind_timing_i(data_ind_timing),
    .data_ind_timing_i_t0(data_ind_timing_t0),
    .div_en_i(div_en_ex),
    .div_en_i_t0(div_en_ex_t0),
    .div_sel_i(div_sel_ex),
    .div_sel_i_t0(div_sel_ex_t0),
    .ex_valid_o(ex_valid),
    .ex_valid_o_t0(ex_valid_t0),
    .imd_val_d_o(imd_val_d_ex),
    .imd_val_d_o_t0(imd_val_d_ex_t0),
    .imd_val_q_i(imd_val_q_ex),
    .imd_val_q_i_t0(imd_val_q_ex_t0),
    .imd_val_we_o(imd_val_we_ex),
    .imd_val_we_o_t0(imd_val_we_ex_t0),
    .mult_en_i(mult_en_ex),
    .mult_en_i_t0(mult_en_ex_t0),
    .mult_sel_i(mult_sel_ex),
    .mult_sel_i_t0(mult_sel_ex_t0),
    .multdiv_operand_a_i(multdiv_operand_a_ex),
    .multdiv_operand_a_i_t0(multdiv_operand_a_ex_t0),
    .multdiv_operand_b_i(multdiv_operand_b_ex),
    .multdiv_operand_b_i_t0(multdiv_operand_b_ex_t0),
    .multdiv_operator_i(multdiv_operator_ex),
    .multdiv_operator_i_t0(multdiv_operator_ex_t0),
    .multdiv_ready_id_i(multdiv_ready_id),
    .multdiv_ready_id_i_t0(multdiv_ready_id_t0),
    .multdiv_signed_mode_i(multdiv_signed_mode_ex),
    .multdiv_signed_mode_i_t0(multdiv_signed_mode_ex_t0),
    .result_ex_o(result_ex),
    .result_ex_o_t0(result_ex_t0),
    .rst_ni(rst_ni)
  );
  paramode8ca0c7d43bf57ed8b25d9c329a7f7eeb115685cauxy_ibex_id_stage  id_stage_i (
    .alu_operand_a_ex_o(alu_operand_a_ex),
    .alu_operand_a_ex_o_t0(alu_operand_a_ex_t0),
    .alu_operand_b_ex_o(alu_operand_b_ex),
    .alu_operand_b_ex_o_t0(alu_operand_b_ex_t0),
    .alu_operator_ex_o(alu_operator_ex),
    .alu_operator_ex_o_t0(alu_operator_ex_t0),
    .branch_decision_i(branch_decision),
    .branch_decision_i_t0(branch_decision_t0),
    .bt_a_operand_o(bt_a_operand),
    .bt_a_operand_o_t0(bt_a_operand_t0),
    .bt_b_operand_o(bt_b_operand),
    .bt_b_operand_o_t0(bt_b_operand_t0),
    .clk_i(clk_i),
    .csr_access_o(csr_access),
    .csr_access_o_t0(csr_access_t0),
    .csr_mstatus_mie_i(csr_mstatus_mie),
    .csr_mstatus_mie_i_t0(csr_mstatus_mie_t0),
    .csr_mstatus_tw_i(csr_mstatus_tw),
    .csr_mstatus_tw_i_t0(csr_mstatus_tw_t0),
    .csr_mtval_o(csr_mtval),
    .csr_mtval_o_t0(csr_mtval_t0),
    .csr_op_en_o(csr_op_en),
    .csr_op_en_o_t0(csr_op_en_t0),
    .csr_op_o(csr_op),
    .csr_op_o_t0(csr_op_t0),
    .csr_rdata_i(csr_rdata),
    .csr_rdata_i_t0(csr_rdata_t0),
    .csr_restore_dret_id_o(csr_restore_dret_id),
    .csr_restore_dret_id_o_t0(csr_restore_dret_id_t0),
    .csr_restore_mret_id_o(csr_restore_mret_id),
    .csr_restore_mret_id_o_t0(csr_restore_mret_id_t0),
    .csr_save_cause_o(csr_save_cause),
    .csr_save_cause_o_t0(csr_save_cause_t0),
    .csr_save_id_o(csr_save_id),
    .csr_save_id_o_t0(csr_save_id_t0),
    .csr_save_if_o(csr_save_if),
    .csr_save_if_o_t0(csr_save_if_t0),
    .csr_save_wb_o(csr_save_wb),
    .csr_save_wb_o_t0(csr_save_wb_t0),
    .ctrl_busy_o(ctrl_busy),
    .ctrl_busy_o_t0(ctrl_busy_t0),
    .data_ind_timing_i(data_ind_timing),
    .data_ind_timing_i_t0(data_ind_timing_t0),
    .debug_cause_o(debug_cause),
    .debug_cause_o_t0(debug_cause_t0),
    .debug_csr_save_o(debug_csr_save),
    .debug_csr_save_o_t0(debug_csr_save_t0),
    .debug_ebreakm_i(debug_ebreakm),
    .debug_ebreakm_i_t0(debug_ebreakm_t0),
    .debug_ebreaku_i(debug_ebreaku),
    .debug_ebreaku_i_t0(debug_ebreaku_t0),
    .debug_mode_o(debug_mode),
    .debug_mode_o_t0(debug_mode_t0),
    .debug_req_i(debug_req_i),
    .debug_req_i_t0(debug_req_i_t0),
    .debug_single_step_i(debug_single_step),
    .debug_single_step_i_t0(debug_single_step_t0),
    .div_en_ex_o(div_en_ex),
    .div_en_ex_o_t0(div_en_ex_t0),
    .div_sel_ex_o(div_sel_ex),
    .div_sel_ex_o_t0(div_sel_ex_t0),
    .en_wb_o(en_wb),
    .en_wb_o_t0(en_wb_t0),
    .ex_valid_i(ex_valid),
    .ex_valid_i_t0(ex_valid_t0),
    .exc_cause_o(exc_cause),
    .exc_cause_o_t0(exc_cause_t0),
    .exc_pc_mux_o(exc_pc_mux_id),
    .exc_pc_mux_o_t0(exc_pc_mux_id_t0),
    .icache_inval_o(icache_inval),
    .icache_inval_o_t0(icache_inval_t0),
    .id_in_ready_o(id_in_ready),
    .id_in_ready_o_t0(id_in_ready_t0),
    .illegal_c_insn_i(illegal_c_insn_id),
    .illegal_c_insn_i_t0(illegal_c_insn_id_t0),
    .illegal_csr_insn_i(illegal_csr_insn_id),
    .illegal_csr_insn_i_t0(illegal_csr_insn_id_t0),
    .illegal_insn_o(illegal_insn_id),
    .illegal_insn_o_t0(illegal_insn_id_t0),
    .imd_val_d_ex_i(imd_val_d_ex),
    .imd_val_d_ex_i_t0(imd_val_d_ex_t0),
    .imd_val_q_ex_o(imd_val_q_ex),
    .imd_val_q_ex_o_t0(imd_val_q_ex_t0),
    .imd_val_we_ex_i(imd_val_we_ex),
    .imd_val_we_ex_i_t0(imd_val_we_ex_t0),
    .instr_bp_taken_i(instr_bp_taken_id),
    .instr_bp_taken_i_t0(instr_bp_taken_id_t0),
    .instr_fetch_err_i(instr_fetch_err),
    .instr_fetch_err_i_t0(instr_fetch_err_t0),
    .instr_fetch_err_plus2_i(instr_fetch_err_plus2),
    .instr_fetch_err_plus2_i_t0(instr_fetch_err_plus2_t0),
    .instr_first_cycle_id_o(instr_first_cycle_id),
    .instr_first_cycle_id_o_t0(instr_first_cycle_id_t0),
    .instr_id_done_o(instr_id_done),
    .instr_id_done_o_t0(instr_id_done_t0),
    .instr_is_compressed_i(instr_is_compressed_id),
    .instr_is_compressed_i_t0(instr_is_compressed_id_t0),
    .instr_perf_count_id_o(instr_perf_count_id),
    .instr_perf_count_id_o_t0(instr_perf_count_id_t0),
    .instr_rdata_alu_i(instr_rdata_alu_id),
    .instr_rdata_alu_i_t0(instr_rdata_alu_id_t0),
    .instr_rdata_c_i(instr_rdata_c_id),
    .instr_rdata_c_i_t0(instr_rdata_c_id_t0),
    .instr_rdata_i(instr_rdata_id),
    .instr_rdata_i_t0(instr_rdata_id_t0),
    .instr_req_o(instr_req_int),
    .instr_req_o_t0(instr_req_int_t0),
    .instr_type_wb_o(instr_type_wb),
    .instr_type_wb_o_t0(instr_type_wb_t0),
    .instr_valid_clear_o(instr_valid_clear),
    .instr_valid_clear_o_t0(instr_valid_clear_t0),
    .instr_valid_i(instr_valid_id),
    .instr_valid_i_t0(instr_valid_id_t0),
    .irq_nm_i(irq_nm_i),
    .irq_nm_i_t0(irq_nm_i_t0),
    .irq_pending_i(irq_pending_o),
    .irq_pending_i_t0(irq_pending_o_t0),
    .irqs_i(irqs),
    .irqs_i_t0(irqs_t0),
    .lsu_addr_incr_req_i(lsu_addr_incr_req),
    .lsu_addr_incr_req_i_t0(lsu_addr_incr_req_t0),
    .lsu_addr_last_i(lsu_addr_last),
    .lsu_addr_last_i_t0(lsu_addr_last_t0),
    .lsu_load_err_i(lsu_load_err),
    .lsu_load_err_i_t0(lsu_load_err_t0),
    .lsu_req_done_i(lsu_req_done),
    .lsu_req_done_i_t0(lsu_req_done_t0),
    .lsu_req_o(lsu_req),
    .lsu_req_o_t0(lsu_req_t0),
    .lsu_resp_valid_i(lsu_resp_valid),
    .lsu_resp_valid_i_t0(lsu_resp_valid_t0),
    .lsu_sign_ext_o(lsu_sign_ext),
    .lsu_sign_ext_o_t0(lsu_sign_ext_t0),
    .lsu_store_err_i(lsu_store_err),
    .lsu_store_err_i_t0(lsu_store_err_t0),
    .lsu_type_o(lsu_type),
    .lsu_type_o_t0(lsu_type_t0),
    .lsu_wdata_o(lsu_wdata),
    .lsu_wdata_o_t0(lsu_wdata_t0),
    .lsu_we_o(lsu_we),
    .lsu_we_o_t0(lsu_we_t0),
    .mult_en_ex_o(mult_en_ex),
    .mult_en_ex_o_t0(mult_en_ex_t0),
    .mult_sel_ex_o(mult_sel_ex),
    .mult_sel_ex_o_t0(mult_sel_ex_t0),
    .multdiv_operand_a_ex_o(multdiv_operand_a_ex),
    .multdiv_operand_a_ex_o_t0(multdiv_operand_a_ex_t0),
    .multdiv_operand_b_ex_o(multdiv_operand_b_ex),
    .multdiv_operand_b_ex_o_t0(multdiv_operand_b_ex_t0),
    .multdiv_operator_ex_o(multdiv_operator_ex),
    .multdiv_operator_ex_o_t0(multdiv_operator_ex_t0),
    .multdiv_ready_id_o(multdiv_ready_id),
    .multdiv_ready_id_o_t0(multdiv_ready_id_t0),
    .multdiv_signed_mode_ex_o(multdiv_signed_mode_ex),
    .multdiv_signed_mode_ex_o_t0(multdiv_signed_mode_ex_t0),
    .nmi_mode_o(nmi_mode),
    .nmi_mode_o_t0(nmi_mode_t0),
    .nt_branch_mispredict_o(nt_branch_mispredict),
    .nt_branch_mispredict_o_t0(nt_branch_mispredict_t0),
    .outstanding_load_wb_i(outstanding_load_wb),
    .outstanding_load_wb_i_t0(outstanding_load_wb_t0),
    .outstanding_store_wb_i(outstanding_store_wb),
    .outstanding_store_wb_i_t0(outstanding_store_wb_t0),
    .pc_id_i(pc_id),
    .pc_id_i_t0(pc_id_t0),
    .pc_mux_o(pc_mux_id),
    .pc_mux_o_t0(pc_mux_id_t0),
    .pc_set_o(pc_set),
    .pc_set_o_t0(pc_set_t0),
    .pc_set_spec_o(pc_set_spec),
    .pc_set_spec_o_t0(pc_set_spec_t0),
    .perf_branch_o(perf_branch),
    .perf_branch_o_t0(perf_branch_t0),
    .perf_div_wait_o(perf_div_wait),
    .perf_div_wait_o_t0(perf_div_wait_t0),
    .perf_dside_wait_o(perf_dside_wait),
    .perf_dside_wait_o_t0(perf_dside_wait_t0),
    .perf_jump_o(perf_jump),
    .perf_jump_o_t0(perf_jump_t0),
    .perf_mul_wait_o(perf_mul_wait),
    .perf_mul_wait_o_t0(perf_mul_wait_t0),
    .perf_tbranch_o(perf_tbranch),
    .perf_tbranch_o_t0(perf_tbranch_t0),
    .priv_mode_i(priv_mode_id),
    .priv_mode_i_t0(priv_mode_id_t0),
    .ready_wb_i(ready_wb),
    .ready_wb_i_t0(ready_wb_t0),
    .result_ex_i(result_ex),
    .result_ex_i_t0(result_ex_t0),
    .rf_raddr_a_o(rf_raddr_a_o),
    .rf_raddr_a_o_t0(rf_raddr_a_o_t0),
    .rf_raddr_b_o(rf_raddr_b_o),
    .rf_raddr_b_o_t0(rf_raddr_b_o_t0),
    .rf_rd_a_wb_match_o(\gen_no_regfile_ecc.unused_rf_rd_a_wb_match ),
    .rf_rd_a_wb_match_o_t0(\gen_no_regfile_ecc.unused_rf_rd_a_wb_match_t0 ),
    .rf_rd_b_wb_match_o(\gen_no_regfile_ecc.unused_rf_rd_b_wb_match ),
    .rf_rd_b_wb_match_o_t0(\gen_no_regfile_ecc.unused_rf_rd_b_wb_match_t0 ),
    .rf_rdata_a_i(rf_rdata_a_ecc_i),
    .rf_rdata_a_i_t0(rf_rdata_a_ecc_i_t0),
    .rf_rdata_b_i(rf_rdata_b_ecc_i),
    .rf_rdata_b_i_t0(rf_rdata_b_ecc_i_t0),
    .rf_ren_a_o(\gen_no_regfile_ecc.unused_rf_ren_a ),
    .rf_ren_a_o_t0(\gen_no_regfile_ecc.unused_rf_ren_a_t0 ),
    .rf_ren_b_o(\gen_no_regfile_ecc.unused_rf_ren_b ),
    .rf_ren_b_o_t0(\gen_no_regfile_ecc.unused_rf_ren_b_t0 ),
    .rf_waddr_id_o(rf_waddr_id),
    .rf_waddr_id_o_t0(rf_waddr_id_t0),
    .rf_waddr_wb_i(rf_waddr_wb_o),
    .rf_waddr_wb_i_t0(rf_waddr_wb_o_t0),
    .rf_wdata_fwd_wb_i(rf_wdata_fwd_wb),
    .rf_wdata_fwd_wb_i_t0(rf_wdata_fwd_wb_t0),
    .rf_wdata_id_o(rf_wdata_id),
    .rf_wdata_id_o_t0(rf_wdata_id_t0),
    .rf_we_id_o(rf_we_id),
    .rf_we_id_o_t0(rf_we_id_t0),
    .rf_write_wb_i(rf_write_wb),
    .rf_write_wb_i_t0(rf_write_wb_t0),
    .rst_ni(rst_ni),
    .trigger_match_i(trigger_match),
    .trigger_match_i_t0(trigger_match_t0)
  );
  paramod228b056930db4609081e7d118c0624e476409ccbauxy_ibex_if_stage  if_stage_i (
    .boot_addr_i(boot_addr_i),
    .boot_addr_i_t0(boot_addr_i_t0),
    .branch_target_ex_i(branch_target_ex),
    .branch_target_ex_i_t0(branch_target_ex_t0),
    .clk_i(clk_i),
    .csr_depc_i(csr_depc),
    .csr_depc_i_t0(csr_depc_t0),
    .csr_mepc_i(csr_mepc),
    .csr_mepc_i_t0(csr_mepc_t0),
    .csr_mtvec_i(csr_mtvec),
    .csr_mtvec_i_t0(csr_mtvec_t0),
    .csr_mtvec_init_o(csr_mtvec_init),
    .csr_mtvec_init_o_t0(csr_mtvec_init_t0),
    .dummy_instr_en_i(dummy_instr_en),
    .dummy_instr_en_i_t0(dummy_instr_en_t0),
    .dummy_instr_id_o(dummy_instr_id_o),
    .dummy_instr_id_o_t0(dummy_instr_id_o_t0),
    .dummy_instr_mask_i(dummy_instr_mask),
    .dummy_instr_mask_i_t0(dummy_instr_mask_t0),
    .dummy_instr_seed_en_i(dummy_instr_seed_en),
    .dummy_instr_seed_en_i_t0(dummy_instr_seed_en_t0),
    .dummy_instr_seed_i(dummy_instr_seed),
    .dummy_instr_seed_i_t0(dummy_instr_seed_t0),
    .exc_cause(exc_cause),
    .exc_cause_t0(exc_cause_t0),
    .exc_pc_mux_i(exc_pc_mux_id),
    .exc_pc_mux_i_t0(exc_pc_mux_id_t0),
    .ic_data_addr_o(ic_data_addr_o),
    .ic_data_addr_o_t0(ic_data_addr_o_t0),
    .ic_data_rdata_i(ic_data_rdata_i),
    .ic_data_rdata_i_t0(ic_data_rdata_i_t0),
    .ic_data_req_o(ic_data_req_o),
    .ic_data_req_o_t0(ic_data_req_o_t0),
    .ic_data_wdata_o(ic_data_wdata_o),
    .ic_data_wdata_o_t0(ic_data_wdata_o_t0),
    .ic_data_write_o(ic_data_write_o),
    .ic_data_write_o_t0(ic_data_write_o_t0),
    .ic_tag_addr_o(ic_tag_addr_o),
    .ic_tag_addr_o_t0(ic_tag_addr_o_t0),
    .ic_tag_rdata_i(ic_tag_rdata_i),
    .ic_tag_rdata_i_t0(ic_tag_rdata_i_t0),
    .ic_tag_req_o(ic_tag_req_o),
    .ic_tag_req_o_t0(ic_tag_req_o_t0),
    .ic_tag_wdata_o(ic_tag_wdata_o),
    .ic_tag_wdata_o_t0(ic_tag_wdata_o_t0),
    .ic_tag_write_o(ic_tag_write_o),
    .ic_tag_write_o_t0(ic_tag_write_o_t0),
    .icache_enable_i(icache_enable),
    .icache_enable_i_t0(icache_enable_t0),
    .icache_inval_i(icache_inval),
    .icache_inval_i_t0(icache_inval_t0),
    .id_in_ready_i(id_in_ready),
    .id_in_ready_i_t0(id_in_ready_t0),
    .if_busy_o(if_busy),
    .if_busy_o_t0(if_busy_t0),
    .illegal_c_insn_id_o(illegal_c_insn_id),
    .illegal_c_insn_id_o_t0(illegal_c_insn_id_t0),
    .instr_addr_o(instr_addr_o),
    .instr_addr_o_t0(instr_addr_o_t0),
    .instr_bp_taken_o(instr_bp_taken_id),
    .instr_bp_taken_o_t0(instr_bp_taken_id_t0),
    .instr_err_i(instr_err_i),
    .instr_err_i_t0(instr_err_i_t0),
    .instr_fetch_err_o(instr_fetch_err),
    .instr_fetch_err_o_t0(instr_fetch_err_t0),
    .instr_fetch_err_plus2_o(instr_fetch_err_plus2),
    .instr_fetch_err_plus2_o_t0(instr_fetch_err_plus2_t0),
    .instr_gnt_i(instr_gnt_i),
    .instr_gnt_i_t0(instr_gnt_i_t0),
    .instr_is_compressed_id_o(instr_is_compressed_id),
    .instr_is_compressed_id_o_t0(instr_is_compressed_id_t0),
    .instr_new_id_o(instr_new_id),
    .instr_new_id_o_t0(instr_new_id_t0),
    .instr_pmp_err_i(1'h0),
    .instr_pmp_err_i_t0(1'h0),
    .instr_rdata_alu_id_o(instr_rdata_alu_id),
    .instr_rdata_alu_id_o_t0(instr_rdata_alu_id_t0),
    .instr_rdata_c_id_o(instr_rdata_c_id),
    .instr_rdata_c_id_o_t0(instr_rdata_c_id_t0),
    .instr_rdata_i(instr_rdata_i),
    .instr_rdata_i_t0(instr_rdata_i_t0),
    .instr_rdata_id_o(instr_rdata_id),
    .instr_rdata_id_o_t0(instr_rdata_id_t0),
    .instr_req_o(instr_req_o),
    .instr_req_o_t0(instr_req_o_t0),
    .instr_rvalid_i(instr_rvalid_i),
    .instr_rvalid_i_t0(instr_rvalid_i_t0),
    .instr_valid_clear_i(instr_valid_clear),
    .instr_valid_clear_i_t0(instr_valid_clear_t0),
    .instr_valid_id_o(instr_valid_id),
    .instr_valid_id_o_t0(instr_valid_id_t0),
    .nt_branch_mispredict_i(nt_branch_mispredict),
    .nt_branch_mispredict_i_t0(nt_branch_mispredict_t0),
    .pc_id_o(pc_id),
    .pc_id_o_t0(pc_id_t0),
    .pc_if_o(pc_if),
    .pc_if_o_t0(pc_if_t0),
    .pc_mismatch_alert_o(pc_mismatch_alert),
    .pc_mismatch_alert_o_t0(pc_mismatch_alert_t0),
    .pc_mux_i(pc_mux_id),
    .pc_mux_i_t0(pc_mux_id_t0),
    .pc_set_i(pc_set),
    .pc_set_i_t0(pc_set_t0),
    .pc_set_spec_i(pc_set_spec),
    .pc_set_spec_i_t0(pc_set_spec_t0),
    .req_i(instr_req_int),
    .req_i_t0(instr_req_int_t0),
    .rst_ni(rst_ni)
  );
  auxy_ibex_load_store_unit load_store_unit_i (
    .adder_result_ex_i(alu_adder_result_ex),
    .adder_result_ex_i_t0(alu_adder_result_ex_t0),
    .addr_incr_req_o(lsu_addr_incr_req),
    .addr_incr_req_o_t0(lsu_addr_incr_req_t0),
    .addr_last_o(lsu_addr_last),
    .addr_last_o_t0(lsu_addr_last_t0),
    .busy_o(lsu_busy),
    .busy_o_t0(lsu_busy_t0),
    .clk_i(clk_i),
    .data_addr_o(data_addr_o),
    .data_addr_o_t0(data_addr_o_t0),
    .data_be_o(data_be_o),
    .data_be_o_t0(data_be_o_t0),
    .data_err_i(data_err_i),
    .data_err_i_t0(data_err_i_t0),
    .data_gnt_i(data_gnt_i),
    .data_gnt_i_t0(data_gnt_i_t0),
    .data_pmp_err_i(1'h0),
    .data_pmp_err_i_t0(1'h0),
    .data_rdata_i(data_rdata_i),
    .data_rdata_i_t0(data_rdata_i_t0),
    .data_req_o(data_req_o),
    .data_req_o_t0(data_req_o_t0),
    .data_rvalid_i(data_rvalid_i),
    .data_rvalid_i_t0(data_rvalid_i_t0),
    .data_wdata_o(data_wdata_o),
    .data_wdata_o_t0(data_wdata_o_t0),
    .data_we_o(data_we_o),
    .data_we_o_t0(data_we_o_t0),
    .load_err_o(lsu_load_err),
    .load_err_o_t0(lsu_load_err_t0),
    .lsu_rdata_o(rf_wdata_lsu),
    .lsu_rdata_o_t0(rf_wdata_lsu_t0),
    .lsu_rdata_valid_o(rf_we_lsu),
    .lsu_rdata_valid_o_t0(rf_we_lsu_t0),
    .lsu_req_done_o(lsu_req_done),
    .lsu_req_done_o_t0(lsu_req_done_t0),
    .lsu_req_i(lsu_req),
    .lsu_req_i_t0(lsu_req_t0),
    .lsu_resp_valid_o(lsu_resp_valid),
    .lsu_resp_valid_o_t0(lsu_resp_valid_t0),
    .lsu_sign_ext_i(lsu_sign_ext),
    .lsu_sign_ext_i_t0(lsu_sign_ext_t0),
    .lsu_type_i(lsu_type),
    .lsu_type_i_t0(lsu_type_t0),
    .lsu_wdata_i(lsu_wdata),
    .lsu_wdata_i_t0(lsu_wdata_t0),
    .lsu_we_i(lsu_we),
    .lsu_we_i_t0(lsu_we_t0),
    .perf_load_o(perf_load),
    .perf_load_o_t0(perf_load_t0),
    .perf_store_o(perf_store),
    .perf_store_o_t0(perf_store_t0),
    .rst_ni(rst_ni),
    .store_err_o(lsu_store_err),
    .store_err_o_t0(lsu_store_err_t0)
  );
  paramodauxy_ibex_wb_stageWritebackStage11  wb_stage_i (
    .clk_i(clk_i),
    .en_wb_i(en_wb),
    .en_wb_i_t0(en_wb_t0),
    .instr_done_wb_o(instr_done_wb),
    .instr_done_wb_o_t0(instr_done_wb_t0),
    .instr_is_compressed_id_i(instr_is_compressed_id),
    .instr_is_compressed_id_i_t0(instr_is_compressed_id_t0),
    .instr_perf_count_id_i(instr_perf_count_id),
    .instr_perf_count_id_i_t0(instr_perf_count_id_t0),
    .instr_type_wb_i(instr_type_wb),
    .instr_type_wb_i_t0(instr_type_wb_t0),
    .lsu_resp_err_i(lsu_resp_err),
    .lsu_resp_err_i_t0(lsu_resp_err_t0),
    .lsu_resp_valid_i(lsu_resp_valid),
    .lsu_resp_valid_i_t0(lsu_resp_valid_t0),
    .outstanding_load_wb_o(outstanding_load_wb),
    .outstanding_load_wb_o_t0(outstanding_load_wb_t0),
    .outstanding_store_wb_o(outstanding_store_wb),
    .outstanding_store_wb_o_t0(outstanding_store_wb_t0),
    .pc_id_i(pc_id),
    .pc_id_i_t0(pc_id_t0),
    .pc_wb_o(pc_wb),
    .pc_wb_o_t0(pc_wb_t0),
    .perf_instr_ret_compressed_wb_o(perf_instr_ret_compressed_wb),
    .perf_instr_ret_compressed_wb_o_t0(perf_instr_ret_compressed_wb_t0),
    .perf_instr_ret_wb_o(perf_instr_ret_wb),
    .perf_instr_ret_wb_o_t0(perf_instr_ret_wb_t0),
    .ready_wb_o(ready_wb),
    .ready_wb_o_t0(ready_wb_t0),
    .rf_waddr_id_i(rf_waddr_id),
    .rf_waddr_id_i_t0(rf_waddr_id_t0),
    .rf_waddr_wb_o(rf_waddr_wb_o),
    .rf_waddr_wb_o_t0(rf_waddr_wb_o_t0),
    .rf_wdata_fwd_wb_o(rf_wdata_fwd_wb),
    .rf_wdata_fwd_wb_o_t0(rf_wdata_fwd_wb_t0),
    .rf_wdata_id_i(rf_wdata_id),
    .rf_wdata_id_i_t0(rf_wdata_id_t0),
    .rf_wdata_lsu_i(rf_wdata_lsu),
    .rf_wdata_lsu_i_t0(rf_wdata_lsu_t0),
    .rf_wdata_wb_o(rf_wdata_wb_ecc_o),
    .rf_wdata_wb_o_t0(rf_wdata_wb_ecc_o_t0),
    .rf_we_id_i(rf_we_id),
    .rf_we_id_i_t0(rf_we_id_t0),
    .rf_we_lsu_i(rf_we_lsu),
    .rf_we_lsu_i_t0(rf_we_lsu_t0),
    .rf_we_wb_o(rf_we_wb_o),
    .rf_we_wb_o_t0(rf_we_wb_o_t0),
    .rf_write_wb_o(rf_write_wb),
    .rf_write_wb_o_t0(rf_write_wb_t0),
    .rst_ni(rst_ni)
  );
  assign alert_minor_o = 1'h0;
  assign alert_minor_o_t0 = 1'h0;
  assign crash_dump_o = { pc_id, pc_if, lsu_addr_last, csr_mepc };
  assign crash_dump_o_t0 = { pc_id_t0, pc_if_t0, lsu_addr_last_t0, csr_mepc_t0 };
endmodule

module paramod16bd66fd1d1dbd7c4dd1efdb08bf1560b5c5007aauxy_ibex_register_file_ff (clk_i, rst_ni, test_en_i, dummy_instr_id_i, raddr_a_i, rdata_a_o, raddr_b_i, rdata_b_o, waddr_a_i, wdata_a_i, we_a_i, we_a_i_t0, wdata_a_i_t0, waddr_a_i_t0, test_en_i_t0, rdata_b_o_t0, rdata_a_o_t0, raddr_b_i_t0, raddr_a_i_t0, dummy_instr_id_i_t0);
  wire _0000_;
  wire _0001_;
  wire _0002_;
  wire _0003_;
  wire _0004_;
  wire _0005_;
  wire _0006_;
  wire _0007_;
  wire _0008_;
  wire _0009_;
  wire _0010_;
  wire _0011_;
  wire _0012_;
  wire _0013_;
  wire _0014_;
  wire _0015_;
  wire _0016_;
  wire _0017_;
  wire _0018_;
  wire _0019_;
  wire _0020_;
  wire _0021_;
  wire _0022_;
  wire _0023_;
  wire _0024_;
  wire _0025_;
  wire _0026_;
  wire _0027_;
  wire _0028_;
  wire _0029_;
  wire _0030_;
  wire [4:0] _0031_;
  wire _0032_;
  wire _0033_;
  wire _0034_;
  wire [31:0] _0035_;
  wire [31:0] _0036_;
  wire [31:0] _0037_;
  wire [31:0] _0038_;
  wire [31:0] _0039_;
  wire [31:0] _0040_;
  wire [31:0] _0041_;
  wire [31:0] _0042_;
  wire [31:0] _0043_;
  wire [31:0] _0044_;
  wire [31:0] _0045_;
  wire [31:0] _0046_;
  wire [31:0] _0047_;
  wire [31:0] _0048_;
  wire [31:0] _0049_;
  wire [31:0] _0050_;
  wire [31:0] _0051_;
  wire [31:0] _0052_;
  wire [31:0] _0053_;
  wire [31:0] _0054_;
  wire [31:0] _0055_;
  wire [31:0] _0056_;
  wire [31:0] _0057_;
  wire [31:0] _0058_;
  wire [31:0] _0059_;
  wire [31:0] _0060_;
  wire [31:0] _0061_;
  wire [31:0] _0062_;
  wire [31:0] _0063_;
  wire [31:0] _0064_;
  wire [31:0] _0065_;
  wire [31:0] _0066_;
  wire [31:0] _0067_;
  wire [31:0] _0068_;
  wire [31:0] _0069_;
  wire [31:0] _0070_;
  wire [31:0] _0071_;
  wire [31:0] _0072_;
  wire [31:0] _0073_;
  wire [31:0] _0074_;
  wire [31:0] _0075_;
  wire [31:0] _0076_;
  wire [31:0] _0077_;
  wire [31:0] _0078_;
  wire [31:0] _0079_;
  wire [31:0] _0080_;
  wire [31:0] _0081_;
  wire [31:0] _0082_;
  wire [31:0] _0083_;
  wire [31:0] _0084_;
  wire [31:0] _0085_;
  wire [31:0] _0086_;
  wire [31:0] _0087_;
  wire [31:0] _0088_;
  wire [31:0] _0089_;
  wire [31:0] _0090_;
  wire [31:0] _0091_;
  wire [31:0] _0092_;
  wire [31:0] _0093_;
  wire [31:0] _0094_;
  wire [31:0] _0095_;
  wire [31:0] _0096_;
  wire [31:0] _0097_;
  wire [31:0] _0098_;
  wire [31:0] _0099_;
  wire [31:0] _0100_;
  wire [31:0] _0101_;
  wire [31:0] _0102_;
  wire [31:0] _0103_;
  wire [31:0] _0104_;
  wire [31:0] _0105_;
  wire [31:0] _0106_;
  wire [31:0] _0107_;
  wire [31:0] _0108_;
  wire [31:0] _0109_;
  wire [31:0] _0110_;
  wire [31:0] _0111_;
  wire [31:0] _0112_;
  wire [31:0] _0113_;
  wire [31:0] _0114_;
  wire [31:0] _0115_;
  wire [31:0] _0116_;
  wire [31:0] _0117_;
  wire [31:0] _0118_;
  wire [31:0] _0119_;
  wire [31:0] _0120_;
  wire [31:0] _0121_;
  wire [31:0] _0122_;
  wire [31:0] _0123_;
  wire [31:0] _0124_;
  wire [31:0] _0125_;
  wire [31:0] _0126_;
  wire [31:0] _0127_;
  wire [4:0] _0128_;
  wire [4:0] _0129_;
  wire [4:0] _0130_;
  wire [4:0] _0131_;
  wire [4:0] _0132_;
  wire [4:0] _0133_;
  wire [4:0] _0134_;
  wire [4:0] _0135_;
  wire [4:0] _0136_;
  wire [4:0] _0137_;
  wire [4:0] _0138_;
  wire [4:0] _0139_;
  wire [4:0] _0140_;
  wire [4:0] _0141_;
  wire [4:0] _0142_;
  wire [4:0] _0143_;
  wire [4:0] _0144_;
  wire [4:0] _0145_;
  wire [4:0] _0146_;
  wire [4:0] _0147_;
  wire [4:0] _0148_;
  wire [4:0] _0149_;
  wire [4:0] _0150_;
  wire [4:0] _0151_;
  wire [4:0] _0152_;
  wire [4:0] _0153_;
  wire [4:0] _0154_;
  wire [4:0] _0155_;
  wire [4:0] _0156_;
  wire [4:0] _0157_;
  wire [4:0] _0158_;
  wire [4:0] _0159_;
  wire _0160_;
  wire _0161_;
  wire _0162_;
  wire _0163_;
  wire _0164_;
  wire _0165_;
  wire _0166_;
  wire _0167_;
  wire _0168_;
  wire _0169_;
  wire _0170_;
  wire _0171_;
  wire _0172_;
  wire _0173_;
  wire _0174_;
  wire _0175_;
  wire _0176_;
  wire _0177_;
  wire _0178_;
  wire _0179_;
  wire _0180_;
  wire _0181_;
  wire _0182_;
  wire _0183_;
  wire _0184_;
  wire _0185_;
  wire _0186_;
  wire _0187_;
  wire _0188_;
  wire _0189_;
  wire _0190_;
  wire _0191_;
  wire _0192_;
  wire _0193_;
  wire _0194_;
  wire _0195_;
  wire _0196_;
  wire _0197_;
  wire _0198_;
  wire _0199_;
  wire _0200_;
  wire _0201_;
  wire _0202_;
  wire _0203_;
  wire _0204_;
  wire _0205_;
  wire _0206_;
  wire _0207_;
  wire _0208_;
  wire _0209_;
  wire _0210_;
  wire _0211_;
  wire _0212_;
  wire _0213_;
  wire _0214_;
  wire _0215_;
  wire _0216_;
  wire _0217_;
  wire _0218_;
  wire _0219_;
  wire _0220_;
  wire _0221_;
  wire [31:0] _0222_;
  wire [31:0] _0223_;
  wire [31:0] _0224_;
  wire [31:0] _0225_;
  wire [31:0] _0226_;
  wire [31:0] _0227_;
  wire [31:0] _0228_;
  wire [31:0] _0229_;
  wire [31:0] _0230_;
  wire [31:0] _0231_;
  wire [31:0] _0232_;
  wire [31:0] _0233_;
  wire [31:0] _0234_;
  wire [31:0] _0235_;
  wire [31:0] _0236_;
  wire [31:0] _0237_;
  wire [31:0] _0238_;
  wire [31:0] _0239_;
  wire [31:0] _0240_;
  wire [31:0] _0241_;
  wire [31:0] _0242_;
  wire [31:0] _0243_;
  wire [31:0] _0244_;
  wire [31:0] _0245_;
  wire [31:0] _0246_;
  wire [31:0] _0247_;
  wire [31:0] _0248_;
  wire [31:0] _0249_;
  wire [31:0] _0250_;
  wire [31:0] _0251_;
  wire [31:0] _0252_;
  wire [31:0] _0253_;
  wire [31:0] _0254_;
  wire [31:0] _0255_;
  wire [31:0] _0256_;
  wire [31:0] _0257_;
  wire [31:0] _0258_;
  wire [31:0] _0259_;
  wire [31:0] _0260_;
  wire [31:0] _0261_;
  wire [31:0] _0262_;
  wire [31:0] _0263_;
  wire [31:0] _0264_;
  wire [31:0] _0265_;
  wire [31:0] _0266_;
  wire [31:0] _0267_;
  wire [31:0] _0268_;
  wire [31:0] _0269_;
  wire [31:0] _0270_;
  wire [31:0] _0271_;
  wire [31:0] _0272_;
  wire [31:0] _0273_;
  wire [31:0] _0274_;
  wire [31:0] _0275_;
  wire [31:0] _0276_;
  wire [31:0] _0277_;
  wire [31:0] _0278_;
  wire [31:0] _0279_;
  wire [31:0] _0280_;
  wire [31:0] _0281_;
  wire [31:0] _0282_;
  wire [31:0] _0283_;
  wire [31:0] _0284_;
  wire [31:0] _0285_;
  wire [31:0] _0286_;
  wire [31:0] _0287_;
  wire [31:0] _0288_;
  wire [31:0] _0289_;
  wire [31:0] _0290_;
  wire [31:0] _0291_;
  wire [31:0] _0292_;
  wire [31:0] _0293_;
  wire [31:0] _0294_;
  wire [31:0] _0295_;
  wire [31:0] _0296_;
  wire [31:0] _0297_;
  wire [31:0] _0298_;
  wire [31:0] _0299_;
  wire [31:0] _0300_;
  wire [31:0] _0301_;
  wire [31:0] _0302_;
  wire [31:0] _0303_;
  wire [31:0] _0304_;
  wire [31:0] _0305_;
  wire [31:0] _0306_;
  wire [31:0] _0307_;
  wire [31:0] _0308_;
  wire [31:0] _0309_;
  wire [31:0] _0310_;
  wire [31:0] _0311_;
  wire [31:0] _0312_;
  wire [31:0] _0313_;
  wire [31:0] _0314_;
  wire [31:0] _0315_;
  wire [31:0] _0316_;
  wire [31:0] _0317_;
  wire [31:0] _0318_;
  wire [31:0] _0319_;
  wire [31:0] _0320_;
  wire [31:0] _0321_;
  wire [31:0] _0322_;
  wire [31:0] _0323_;
  wire [31:0] _0324_;
  wire [31:0] _0325_;
  wire [31:0] _0326_;
  wire [31:0] _0327_;
  wire [31:0] _0328_;
  wire [31:0] _0329_;
  wire [31:0] _0330_;
  wire [31:0] _0331_;
  wire [31:0] _0332_;
  wire [31:0] _0333_;
  wire [31:0] _0334_;
  wire [31:0] _0335_;
  wire [31:0] _0336_;
  wire [31:0] _0337_;
  wire [31:0] _0338_;
  wire [31:0] _0339_;
  wire [31:0] _0340_;
  wire [31:0] _0341_;
  wire [31:0] _0342_;
  wire [31:0] _0343_;
  wire [31:0] _0344_;
  wire [31:0] _0345_;
  wire _0346_;
  wire _0347_;
  wire _0348_;
  wire _0349_;
  wire _0350_;
  wire _0351_;
  wire _0352_;
  wire _0353_;
  wire _0354_;
  wire _0355_;
  wire _0356_;
  wire _0357_;
  wire _0358_;
  wire _0359_;
  wire _0360_;
  wire _0361_;
  wire _0362_;
  wire _0363_;
  wire _0364_;
  wire _0365_;
  wire _0366_;
  wire _0367_;
  wire _0368_;
  wire _0369_;
  wire _0370_;
  wire _0371_;
  wire _0372_;
  wire _0373_;
  wire _0374_;
  wire _0375_;
  wire _0376_;
  wire [31:0] _0377_;
  wire [31:0] _0378_;
  wire [31:0] _0379_;
  wire [31:0] _0380_;
  wire [31:0] _0381_;
  wire [31:0] _0382_;
  wire [31:0] _0383_;
  wire [31:0] _0384_;
  wire [31:0] _0385_;
  wire [31:0] _0386_;
  wire [31:0] _0387_;
  wire [31:0] _0388_;
  wire [31:0] _0389_;
  wire [31:0] _0390_;
  wire [31:0] _0391_;
  wire [31:0] _0392_;
  wire [31:0] _0393_;
  wire [31:0] _0394_;
  wire [31:0] _0395_;
  wire [31:0] _0396_;
  wire [31:0] _0397_;
  wire [31:0] _0398_;
  wire [31:0] _0399_;
  wire [31:0] _0400_;
  wire [31:0] _0401_;
  wire [31:0] _0402_;
  wire [31:0] _0403_;
  wire [31:0] _0404_;
  wire [31:0] _0405_;
  wire [31:0] _0406_;
  wire [31:0] _0407_;
  wire _0408_;
  wire _0409_;
  wire _0410_;
  wire _0411_;
  wire _0412_;
  wire _0413_;
  wire _0414_;
  wire _0415_;
  wire _0416_;
  wire _0417_;
  wire _0418_;
  wire _0419_;
  wire _0420_;
  wire _0421_;
  wire _0422_;
  wire _0423_;
  wire _0424_;
  wire _0425_;
  wire _0426_;
  wire _0427_;
  wire _0428_;
  wire _0429_;
  wire _0430_;
  wire _0431_;
  wire _0432_;
  wire _0433_;
  wire _0434_;
  wire _0435_;
  wire _0436_;
  wire _0437_;
  wire _0438_;
  wire [31:0] _0439_;
  wire [31:0] _0440_;
  wire _0441_;
  wire _0442_;
  wire _0443_;
  wire _0444_;
  wire _0445_;
  wire _0446_;
  wire _0447_;
  wire _0448_;
  wire _0449_;
  wire _0450_;
  wire _0451_;
  wire _0452_;
  wire _0453_;
  wire _0454_;
  wire _0455_;
  wire _0456_;
  wire _0457_;
  wire _0458_;
  wire _0459_;
  wire _0460_;
  wire _0461_;
  wire _0462_;
  wire _0463_;
  wire _0464_;
  wire _0465_;
  wire _0466_;
  wire _0467_;
  wire _0468_;
  wire _0469_;
  wire _0470_;
  wire _0471_;
  wire _0472_;
  wire _0473_;
  wire _0474_;
  wire _0475_;
  wire _0476_;
  wire _0477_;
  wire _0478_;
  wire _0479_;
  wire _0480_;
  wire _0481_;
  wire _0482_;
  wire _0483_;
  wire _0484_;
  wire _0485_;
  wire _0486_;
  wire _0487_;
  wire _0488_;
  wire _0489_;
  wire _0490_;
  wire _0491_;
  wire _0492_;
  wire _0493_;
  wire _0494_;
  wire _0495_;
  wire _0496_;
  wire _0497_;
  wire _0498_;
  wire _0499_;
  wire _0500_;
  wire _0501_;
  wire _0502_;
  input clk_i;
  wire clk_i;
  input dummy_instr_id_i;
  wire dummy_instr_id_i;
  input dummy_instr_id_i_t0;
  wire dummy_instr_id_i_t0;
  input [4:0] raddr_a_i;
  wire [4:0] raddr_a_i;
  input [4:0] raddr_a_i_t0;
  wire [4:0] raddr_a_i_t0;
  input [4:0] raddr_b_i;
  wire [4:0] raddr_b_i;
  input [4:0] raddr_b_i_t0;
  wire [4:0] raddr_b_i_t0;
  output [31:0] rdata_a_o;
  wire [31:0] rdata_a_o;
  output [31:0] rdata_a_o_t0;
  wire [31:0] rdata_a_o_t0;
  output [31:0] rdata_b_o;
  wire [31:0] rdata_b_o;
  output [31:0] rdata_b_o_t0;
  wire [31:0] rdata_b_o_t0;
  wire [1023:0] rf_reg;
  wire [1023:0] rf_reg_t0;
  input rst_ni;
  wire rst_ni;
  input test_en_i;
  wire test_en_i;
  input test_en_i_t0;
  wire test_en_i_t0;
  input [4:0] waddr_a_i;
  wire [4:0] waddr_a_i;
  input [4:0] waddr_a_i_t0;
  wire [4:0] waddr_a_i_t0;
  input [31:0] wdata_a_i;
  wire [31:0] wdata_a_i;
  input [31:0] wdata_a_i_t0;
  wire [31:0] wdata_a_i_t0;
  wire [31:1] we_a_dec;
  wire [31:1] we_a_dec_t0;
  input we_a_i;
  wire we_a_i;
  input we_a_i_t0;
  wire we_a_i_t0;
  assign _0000_ = ~ we_a_dec[1];
  assign _0001_ = ~ we_a_dec[2];
  assign _0002_ = ~ we_a_dec[31];
  assign _0003_ = ~ we_a_dec[30];
  assign _0004_ = ~ we_a_dec[29];
  assign _0005_ = ~ we_a_dec[28];
  assign _0006_ = ~ we_a_dec[27];
  assign _0007_ = ~ we_a_dec[26];
  assign _0008_ = ~ we_a_dec[25];
  assign _0009_ = ~ we_a_dec[24];
  assign _0010_ = ~ we_a_dec[23];
  assign _0011_ = ~ we_a_dec[22];
  assign _0012_ = ~ we_a_dec[21];
  assign _0013_ = ~ we_a_dec[20];
  assign _0014_ = ~ we_a_dec[19];
  assign _0015_ = ~ we_a_dec[18];
  assign _0016_ = ~ we_a_dec[17];
  assign _0017_ = ~ we_a_dec[16];
  assign _0018_ = ~ we_a_dec[15];
  assign _0019_ = ~ we_a_dec[14];
  assign _0020_ = ~ we_a_dec[13];
  assign _0021_ = ~ we_a_dec[12];
  assign _0022_ = ~ we_a_dec[11];
  assign _0023_ = ~ we_a_dec[10];
  assign _0024_ = ~ we_a_dec[9];
  assign _0025_ = ~ we_a_dec[8];
  assign _0026_ = ~ we_a_dec[7];
  assign _0027_ = ~ we_a_dec[6];
  assign _0028_ = ~ we_a_dec[5];
  assign _0029_ = ~ we_a_dec[4];
  assign _0030_ = ~ we_a_dec[3];
  assign _0377_ = wdata_a_i ^ rf_reg[63:32];
  assign _0378_ = wdata_a_i ^ rf_reg[95:64];
  assign _0379_ = wdata_a_i ^ rf_reg[1023:992];
  assign _0380_ = wdata_a_i ^ rf_reg[991:960];
  assign _0381_ = wdata_a_i ^ rf_reg[959:928];
  assign _0382_ = wdata_a_i ^ rf_reg[927:896];
  assign _0383_ = wdata_a_i ^ rf_reg[895:864];
  assign _0384_ = wdata_a_i ^ rf_reg[863:832];
  assign _0385_ = wdata_a_i ^ rf_reg[831:800];
  assign _0386_ = wdata_a_i ^ rf_reg[799:768];
  assign _0387_ = wdata_a_i ^ rf_reg[767:736];
  assign _0388_ = wdata_a_i ^ rf_reg[735:704];
  assign _0389_ = wdata_a_i ^ rf_reg[703:672];
  assign _0390_ = wdata_a_i ^ rf_reg[671:640];
  assign _0391_ = wdata_a_i ^ rf_reg[639:608];
  assign _0392_ = wdata_a_i ^ rf_reg[607:576];
  assign _0393_ = wdata_a_i ^ rf_reg[575:544];
  assign _0394_ = wdata_a_i ^ rf_reg[543:512];
  assign _0395_ = wdata_a_i ^ rf_reg[511:480];
  assign _0396_ = wdata_a_i ^ rf_reg[479:448];
  assign _0397_ = wdata_a_i ^ rf_reg[447:416];
  assign _0398_ = wdata_a_i ^ rf_reg[415:384];
  assign _0399_ = wdata_a_i ^ rf_reg[383:352];
  assign _0400_ = wdata_a_i ^ rf_reg[351:320];
  assign _0401_ = wdata_a_i ^ rf_reg[319:288];
  assign _0402_ = wdata_a_i ^ rf_reg[287:256];
  assign _0403_ = wdata_a_i ^ rf_reg[255:224];
  assign _0404_ = wdata_a_i ^ rf_reg[223:192];
  assign _0405_ = wdata_a_i ^ rf_reg[191:160];
  assign _0406_ = wdata_a_i ^ rf_reg[159:128];
  assign _0407_ = wdata_a_i ^ rf_reg[127:96];
  assign _0222_ = wdata_a_i_t0 | rf_reg_t0[63:32];
  assign _0226_ = wdata_a_i_t0 | rf_reg_t0[95:64];
  assign _0230_ = wdata_a_i_t0 | rf_reg_t0[1023:992];
  assign _0234_ = wdata_a_i_t0 | rf_reg_t0[991:960];
  assign _0238_ = wdata_a_i_t0 | rf_reg_t0[959:928];
  assign _0242_ = wdata_a_i_t0 | rf_reg_t0[927:896];
  assign _0246_ = wdata_a_i_t0 | rf_reg_t0[895:864];
  assign _0250_ = wdata_a_i_t0 | rf_reg_t0[863:832];
  assign _0254_ = wdata_a_i_t0 | rf_reg_t0[831:800];
  assign _0258_ = wdata_a_i_t0 | rf_reg_t0[799:768];
  assign _0262_ = wdata_a_i_t0 | rf_reg_t0[767:736];
  assign _0266_ = wdata_a_i_t0 | rf_reg_t0[735:704];
  assign _0270_ = wdata_a_i_t0 | rf_reg_t0[703:672];
  assign _0274_ = wdata_a_i_t0 | rf_reg_t0[671:640];
  assign _0278_ = wdata_a_i_t0 | rf_reg_t0[639:608];
  assign _0282_ = wdata_a_i_t0 | rf_reg_t0[607:576];
  assign _0286_ = wdata_a_i_t0 | rf_reg_t0[575:544];
  assign _0290_ = wdata_a_i_t0 | rf_reg_t0[543:512];
  assign _0294_ = wdata_a_i_t0 | rf_reg_t0[511:480];
  assign _0298_ = wdata_a_i_t0 | rf_reg_t0[479:448];
  assign _0302_ = wdata_a_i_t0 | rf_reg_t0[447:416];
  assign _0306_ = wdata_a_i_t0 | rf_reg_t0[415:384];
  assign _0310_ = wdata_a_i_t0 | rf_reg_t0[383:352];
  assign _0314_ = wdata_a_i_t0 | rf_reg_t0[351:320];
  assign _0318_ = wdata_a_i_t0 | rf_reg_t0[319:288];
  assign _0322_ = wdata_a_i_t0 | rf_reg_t0[287:256];
  assign _0326_ = wdata_a_i_t0 | rf_reg_t0[255:224];
  assign _0330_ = wdata_a_i_t0 | rf_reg_t0[223:192];
  assign _0334_ = wdata_a_i_t0 | rf_reg_t0[191:160];
  assign _0338_ = wdata_a_i_t0 | rf_reg_t0[159:128];
  assign _0342_ = wdata_a_i_t0 | rf_reg_t0[127:96];
  assign _0223_ = _0377_ | _0222_;
  assign _0227_ = _0378_ | _0226_;
  assign _0231_ = _0379_ | _0230_;
  assign _0235_ = _0380_ | _0234_;
  assign _0239_ = _0381_ | _0238_;
  assign _0243_ = _0382_ | _0242_;
  assign _0247_ = _0383_ | _0246_;
  assign _0251_ = _0384_ | _0250_;
  assign _0255_ = _0385_ | _0254_;
  assign _0259_ = _0386_ | _0258_;
  assign _0263_ = _0387_ | _0262_;
  assign _0267_ = _0388_ | _0266_;
  assign _0271_ = _0389_ | _0270_;
  assign _0275_ = _0390_ | _0274_;
  assign _0279_ = _0391_ | _0278_;
  assign _0283_ = _0392_ | _0282_;
  assign _0287_ = _0393_ | _0286_;
  assign _0291_ = _0394_ | _0290_;
  assign _0295_ = _0395_ | _0294_;
  assign _0299_ = _0396_ | _0298_;
  assign _0303_ = _0397_ | _0302_;
  assign _0307_ = _0398_ | _0306_;
  assign _0311_ = _0399_ | _0310_;
  assign _0315_ = _0400_ | _0314_;
  assign _0319_ = _0401_ | _0318_;
  assign _0323_ = _0402_ | _0322_;
  assign _0327_ = _0403_ | _0326_;
  assign _0331_ = _0404_ | _0330_;
  assign _0335_ = _0405_ | _0334_;
  assign _0339_ = _0406_ | _0338_;
  assign _0343_ = _0407_ | _0342_;
  assign _0035_ = { we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1] } & wdata_a_i_t0;
  assign _0038_ = { we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2] } & wdata_a_i_t0;
  assign _0041_ = { we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31] } & wdata_a_i_t0;
  assign _0044_ = { we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30] } & wdata_a_i_t0;
  assign _0047_ = { we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29] } & wdata_a_i_t0;
  assign _0050_ = { we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28] } & wdata_a_i_t0;
  assign _0053_ = { we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27] } & wdata_a_i_t0;
  assign _0056_ = { we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26] } & wdata_a_i_t0;
  assign _0059_ = { we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25] } & wdata_a_i_t0;
  assign _0062_ = { we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24] } & wdata_a_i_t0;
  assign _0065_ = { we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23] } & wdata_a_i_t0;
  assign _0068_ = { we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22] } & wdata_a_i_t0;
  assign _0071_ = { we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21] } & wdata_a_i_t0;
  assign _0074_ = { we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20] } & wdata_a_i_t0;
  assign _0077_ = { we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19] } & wdata_a_i_t0;
  assign _0080_ = { we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18] } & wdata_a_i_t0;
  assign _0083_ = { we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17] } & wdata_a_i_t0;
  assign _0086_ = { we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16] } & wdata_a_i_t0;
  assign _0089_ = { we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15] } & wdata_a_i_t0;
  assign _0092_ = { we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14] } & wdata_a_i_t0;
  assign _0095_ = { we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13] } & wdata_a_i_t0;
  assign _0098_ = { we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12] } & wdata_a_i_t0;
  assign _0101_ = { we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11] } & wdata_a_i_t0;
  assign _0104_ = { we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10] } & wdata_a_i_t0;
  assign _0107_ = { we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9] } & wdata_a_i_t0;
  assign _0110_ = { we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8] } & wdata_a_i_t0;
  assign _0113_ = { we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7] } & wdata_a_i_t0;
  assign _0116_ = { we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6] } & wdata_a_i_t0;
  assign _0119_ = { we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5] } & wdata_a_i_t0;
  assign _0122_ = { we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4] } & wdata_a_i_t0;
  assign _0125_ = { we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3] } & wdata_a_i_t0;
  assign _0036_ = { _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_ } & rf_reg_t0[63:32];
  assign _0039_ = { _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_ } & rf_reg_t0[95:64];
  assign _0042_ = { _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_ } & rf_reg_t0[1023:992];
  assign _0045_ = { _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_ } & rf_reg_t0[991:960];
  assign _0048_ = { _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_ } & rf_reg_t0[959:928];
  assign _0051_ = { _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_ } & rf_reg_t0[927:896];
  assign _0054_ = { _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_ } & rf_reg_t0[895:864];
  assign _0057_ = { _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_ } & rf_reg_t0[863:832];
  assign _0060_ = { _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_ } & rf_reg_t0[831:800];
  assign _0063_ = { _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_ } & rf_reg_t0[799:768];
  assign _0066_ = { _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_ } & rf_reg_t0[767:736];
  assign _0069_ = { _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_ } & rf_reg_t0[735:704];
  assign _0072_ = { _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_ } & rf_reg_t0[703:672];
  assign _0075_ = { _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_ } & rf_reg_t0[671:640];
  assign _0078_ = { _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_ } & rf_reg_t0[639:608];
  assign _0081_ = { _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_ } & rf_reg_t0[607:576];
  assign _0084_ = { _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_ } & rf_reg_t0[575:544];
  assign _0087_ = { _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_ } & rf_reg_t0[543:512];
  assign _0090_ = { _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_ } & rf_reg_t0[511:480];
  assign _0093_ = { _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_ } & rf_reg_t0[479:448];
  assign _0096_ = { _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_ } & rf_reg_t0[447:416];
  assign _0099_ = { _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_ } & rf_reg_t0[415:384];
  assign _0102_ = { _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_ } & rf_reg_t0[383:352];
  assign _0105_ = { _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_ } & rf_reg_t0[351:320];
  assign _0108_ = { _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_ } & rf_reg_t0[319:288];
  assign _0111_ = { _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_ } & rf_reg_t0[287:256];
  assign _0114_ = { _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_ } & rf_reg_t0[255:224];
  assign _0117_ = { _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_ } & rf_reg_t0[223:192];
  assign _0120_ = { _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_ } & rf_reg_t0[191:160];
  assign _0123_ = { _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_ } & rf_reg_t0[159:128];
  assign _0126_ = { _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_ } & rf_reg_t0[127:96];
  assign _0037_ = _0223_ & { we_a_dec_t0[1], we_a_dec_t0[1], we_a_dec_t0[1], we_a_dec_t0[1], we_a_dec_t0[1], we_a_dec_t0[1], we_a_dec_t0[1], we_a_dec_t0[1], we_a_dec_t0[1], we_a_dec_t0[1], we_a_dec_t0[1], we_a_dec_t0[1], we_a_dec_t0[1], we_a_dec_t0[1], we_a_dec_t0[1], we_a_dec_t0[1], we_a_dec_t0[1], we_a_dec_t0[1], we_a_dec_t0[1], we_a_dec_t0[1], we_a_dec_t0[1], we_a_dec_t0[1], we_a_dec_t0[1], we_a_dec_t0[1], we_a_dec_t0[1], we_a_dec_t0[1], we_a_dec_t0[1], we_a_dec_t0[1], we_a_dec_t0[1], we_a_dec_t0[1], we_a_dec_t0[1], we_a_dec_t0[1] };
  assign _0040_ = _0227_ & { we_a_dec_t0[2], we_a_dec_t0[2], we_a_dec_t0[2], we_a_dec_t0[2], we_a_dec_t0[2], we_a_dec_t0[2], we_a_dec_t0[2], we_a_dec_t0[2], we_a_dec_t0[2], we_a_dec_t0[2], we_a_dec_t0[2], we_a_dec_t0[2], we_a_dec_t0[2], we_a_dec_t0[2], we_a_dec_t0[2], we_a_dec_t0[2], we_a_dec_t0[2], we_a_dec_t0[2], we_a_dec_t0[2], we_a_dec_t0[2], we_a_dec_t0[2], we_a_dec_t0[2], we_a_dec_t0[2], we_a_dec_t0[2], we_a_dec_t0[2], we_a_dec_t0[2], we_a_dec_t0[2], we_a_dec_t0[2], we_a_dec_t0[2], we_a_dec_t0[2], we_a_dec_t0[2], we_a_dec_t0[2] };
  assign _0043_ = _0231_ & { we_a_dec_t0[31], we_a_dec_t0[31], we_a_dec_t0[31], we_a_dec_t0[31], we_a_dec_t0[31], we_a_dec_t0[31], we_a_dec_t0[31], we_a_dec_t0[31], we_a_dec_t0[31], we_a_dec_t0[31], we_a_dec_t0[31], we_a_dec_t0[31], we_a_dec_t0[31], we_a_dec_t0[31], we_a_dec_t0[31], we_a_dec_t0[31], we_a_dec_t0[31], we_a_dec_t0[31], we_a_dec_t0[31], we_a_dec_t0[31], we_a_dec_t0[31], we_a_dec_t0[31], we_a_dec_t0[31], we_a_dec_t0[31], we_a_dec_t0[31], we_a_dec_t0[31], we_a_dec_t0[31], we_a_dec_t0[31], we_a_dec_t0[31], we_a_dec_t0[31], we_a_dec_t0[31], we_a_dec_t0[31] };
  assign _0046_ = _0235_ & { we_a_dec_t0[30], we_a_dec_t0[30], we_a_dec_t0[30], we_a_dec_t0[30], we_a_dec_t0[30], we_a_dec_t0[30], we_a_dec_t0[30], we_a_dec_t0[30], we_a_dec_t0[30], we_a_dec_t0[30], we_a_dec_t0[30], we_a_dec_t0[30], we_a_dec_t0[30], we_a_dec_t0[30], we_a_dec_t0[30], we_a_dec_t0[30], we_a_dec_t0[30], we_a_dec_t0[30], we_a_dec_t0[30], we_a_dec_t0[30], we_a_dec_t0[30], we_a_dec_t0[30], we_a_dec_t0[30], we_a_dec_t0[30], we_a_dec_t0[30], we_a_dec_t0[30], we_a_dec_t0[30], we_a_dec_t0[30], we_a_dec_t0[30], we_a_dec_t0[30], we_a_dec_t0[30], we_a_dec_t0[30] };
  assign _0049_ = _0239_ & { we_a_dec_t0[29], we_a_dec_t0[29], we_a_dec_t0[29], we_a_dec_t0[29], we_a_dec_t0[29], we_a_dec_t0[29], we_a_dec_t0[29], we_a_dec_t0[29], we_a_dec_t0[29], we_a_dec_t0[29], we_a_dec_t0[29], we_a_dec_t0[29], we_a_dec_t0[29], we_a_dec_t0[29], we_a_dec_t0[29], we_a_dec_t0[29], we_a_dec_t0[29], we_a_dec_t0[29], we_a_dec_t0[29], we_a_dec_t0[29], we_a_dec_t0[29], we_a_dec_t0[29], we_a_dec_t0[29], we_a_dec_t0[29], we_a_dec_t0[29], we_a_dec_t0[29], we_a_dec_t0[29], we_a_dec_t0[29], we_a_dec_t0[29], we_a_dec_t0[29], we_a_dec_t0[29], we_a_dec_t0[29] };
  assign _0052_ = _0243_ & { we_a_dec_t0[28], we_a_dec_t0[28], we_a_dec_t0[28], we_a_dec_t0[28], we_a_dec_t0[28], we_a_dec_t0[28], we_a_dec_t0[28], we_a_dec_t0[28], we_a_dec_t0[28], we_a_dec_t0[28], we_a_dec_t0[28], we_a_dec_t0[28], we_a_dec_t0[28], we_a_dec_t0[28], we_a_dec_t0[28], we_a_dec_t0[28], we_a_dec_t0[28], we_a_dec_t0[28], we_a_dec_t0[28], we_a_dec_t0[28], we_a_dec_t0[28], we_a_dec_t0[28], we_a_dec_t0[28], we_a_dec_t0[28], we_a_dec_t0[28], we_a_dec_t0[28], we_a_dec_t0[28], we_a_dec_t0[28], we_a_dec_t0[28], we_a_dec_t0[28], we_a_dec_t0[28], we_a_dec_t0[28] };
  assign _0055_ = _0247_ & { we_a_dec_t0[27], we_a_dec_t0[27], we_a_dec_t0[27], we_a_dec_t0[27], we_a_dec_t0[27], we_a_dec_t0[27], we_a_dec_t0[27], we_a_dec_t0[27], we_a_dec_t0[27], we_a_dec_t0[27], we_a_dec_t0[27], we_a_dec_t0[27], we_a_dec_t0[27], we_a_dec_t0[27], we_a_dec_t0[27], we_a_dec_t0[27], we_a_dec_t0[27], we_a_dec_t0[27], we_a_dec_t0[27], we_a_dec_t0[27], we_a_dec_t0[27], we_a_dec_t0[27], we_a_dec_t0[27], we_a_dec_t0[27], we_a_dec_t0[27], we_a_dec_t0[27], we_a_dec_t0[27], we_a_dec_t0[27], we_a_dec_t0[27], we_a_dec_t0[27], we_a_dec_t0[27], we_a_dec_t0[27] };
  assign _0058_ = _0251_ & { we_a_dec_t0[26], we_a_dec_t0[26], we_a_dec_t0[26], we_a_dec_t0[26], we_a_dec_t0[26], we_a_dec_t0[26], we_a_dec_t0[26], we_a_dec_t0[26], we_a_dec_t0[26], we_a_dec_t0[26], we_a_dec_t0[26], we_a_dec_t0[26], we_a_dec_t0[26], we_a_dec_t0[26], we_a_dec_t0[26], we_a_dec_t0[26], we_a_dec_t0[26], we_a_dec_t0[26], we_a_dec_t0[26], we_a_dec_t0[26], we_a_dec_t0[26], we_a_dec_t0[26], we_a_dec_t0[26], we_a_dec_t0[26], we_a_dec_t0[26], we_a_dec_t0[26], we_a_dec_t0[26], we_a_dec_t0[26], we_a_dec_t0[26], we_a_dec_t0[26], we_a_dec_t0[26], we_a_dec_t0[26] };
  assign _0061_ = _0255_ & { we_a_dec_t0[25], we_a_dec_t0[25], we_a_dec_t0[25], we_a_dec_t0[25], we_a_dec_t0[25], we_a_dec_t0[25], we_a_dec_t0[25], we_a_dec_t0[25], we_a_dec_t0[25], we_a_dec_t0[25], we_a_dec_t0[25], we_a_dec_t0[25], we_a_dec_t0[25], we_a_dec_t0[25], we_a_dec_t0[25], we_a_dec_t0[25], we_a_dec_t0[25], we_a_dec_t0[25], we_a_dec_t0[25], we_a_dec_t0[25], we_a_dec_t0[25], we_a_dec_t0[25], we_a_dec_t0[25], we_a_dec_t0[25], we_a_dec_t0[25], we_a_dec_t0[25], we_a_dec_t0[25], we_a_dec_t0[25], we_a_dec_t0[25], we_a_dec_t0[25], we_a_dec_t0[25], we_a_dec_t0[25] };
  assign _0064_ = _0259_ & { we_a_dec_t0[24], we_a_dec_t0[24], we_a_dec_t0[24], we_a_dec_t0[24], we_a_dec_t0[24], we_a_dec_t0[24], we_a_dec_t0[24], we_a_dec_t0[24], we_a_dec_t0[24], we_a_dec_t0[24], we_a_dec_t0[24], we_a_dec_t0[24], we_a_dec_t0[24], we_a_dec_t0[24], we_a_dec_t0[24], we_a_dec_t0[24], we_a_dec_t0[24], we_a_dec_t0[24], we_a_dec_t0[24], we_a_dec_t0[24], we_a_dec_t0[24], we_a_dec_t0[24], we_a_dec_t0[24], we_a_dec_t0[24], we_a_dec_t0[24], we_a_dec_t0[24], we_a_dec_t0[24], we_a_dec_t0[24], we_a_dec_t0[24], we_a_dec_t0[24], we_a_dec_t0[24], we_a_dec_t0[24] };
  assign _0067_ = _0263_ & { we_a_dec_t0[23], we_a_dec_t0[23], we_a_dec_t0[23], we_a_dec_t0[23], we_a_dec_t0[23], we_a_dec_t0[23], we_a_dec_t0[23], we_a_dec_t0[23], we_a_dec_t0[23], we_a_dec_t0[23], we_a_dec_t0[23], we_a_dec_t0[23], we_a_dec_t0[23], we_a_dec_t0[23], we_a_dec_t0[23], we_a_dec_t0[23], we_a_dec_t0[23], we_a_dec_t0[23], we_a_dec_t0[23], we_a_dec_t0[23], we_a_dec_t0[23], we_a_dec_t0[23], we_a_dec_t0[23], we_a_dec_t0[23], we_a_dec_t0[23], we_a_dec_t0[23], we_a_dec_t0[23], we_a_dec_t0[23], we_a_dec_t0[23], we_a_dec_t0[23], we_a_dec_t0[23], we_a_dec_t0[23] };
  assign _0070_ = _0267_ & { we_a_dec_t0[22], we_a_dec_t0[22], we_a_dec_t0[22], we_a_dec_t0[22], we_a_dec_t0[22], we_a_dec_t0[22], we_a_dec_t0[22], we_a_dec_t0[22], we_a_dec_t0[22], we_a_dec_t0[22], we_a_dec_t0[22], we_a_dec_t0[22], we_a_dec_t0[22], we_a_dec_t0[22], we_a_dec_t0[22], we_a_dec_t0[22], we_a_dec_t0[22], we_a_dec_t0[22], we_a_dec_t0[22], we_a_dec_t0[22], we_a_dec_t0[22], we_a_dec_t0[22], we_a_dec_t0[22], we_a_dec_t0[22], we_a_dec_t0[22], we_a_dec_t0[22], we_a_dec_t0[22], we_a_dec_t0[22], we_a_dec_t0[22], we_a_dec_t0[22], we_a_dec_t0[22], we_a_dec_t0[22] };
  assign _0073_ = _0271_ & { we_a_dec_t0[21], we_a_dec_t0[21], we_a_dec_t0[21], we_a_dec_t0[21], we_a_dec_t0[21], we_a_dec_t0[21], we_a_dec_t0[21], we_a_dec_t0[21], we_a_dec_t0[21], we_a_dec_t0[21], we_a_dec_t0[21], we_a_dec_t0[21], we_a_dec_t0[21], we_a_dec_t0[21], we_a_dec_t0[21], we_a_dec_t0[21], we_a_dec_t0[21], we_a_dec_t0[21], we_a_dec_t0[21], we_a_dec_t0[21], we_a_dec_t0[21], we_a_dec_t0[21], we_a_dec_t0[21], we_a_dec_t0[21], we_a_dec_t0[21], we_a_dec_t0[21], we_a_dec_t0[21], we_a_dec_t0[21], we_a_dec_t0[21], we_a_dec_t0[21], we_a_dec_t0[21], we_a_dec_t0[21] };
  assign _0076_ = _0275_ & { we_a_dec_t0[20], we_a_dec_t0[20], we_a_dec_t0[20], we_a_dec_t0[20], we_a_dec_t0[20], we_a_dec_t0[20], we_a_dec_t0[20], we_a_dec_t0[20], we_a_dec_t0[20], we_a_dec_t0[20], we_a_dec_t0[20], we_a_dec_t0[20], we_a_dec_t0[20], we_a_dec_t0[20], we_a_dec_t0[20], we_a_dec_t0[20], we_a_dec_t0[20], we_a_dec_t0[20], we_a_dec_t0[20], we_a_dec_t0[20], we_a_dec_t0[20], we_a_dec_t0[20], we_a_dec_t0[20], we_a_dec_t0[20], we_a_dec_t0[20], we_a_dec_t0[20], we_a_dec_t0[20], we_a_dec_t0[20], we_a_dec_t0[20], we_a_dec_t0[20], we_a_dec_t0[20], we_a_dec_t0[20] };
  assign _0079_ = _0279_ & { we_a_dec_t0[19], we_a_dec_t0[19], we_a_dec_t0[19], we_a_dec_t0[19], we_a_dec_t0[19], we_a_dec_t0[19], we_a_dec_t0[19], we_a_dec_t0[19], we_a_dec_t0[19], we_a_dec_t0[19], we_a_dec_t0[19], we_a_dec_t0[19], we_a_dec_t0[19], we_a_dec_t0[19], we_a_dec_t0[19], we_a_dec_t0[19], we_a_dec_t0[19], we_a_dec_t0[19], we_a_dec_t0[19], we_a_dec_t0[19], we_a_dec_t0[19], we_a_dec_t0[19], we_a_dec_t0[19], we_a_dec_t0[19], we_a_dec_t0[19], we_a_dec_t0[19], we_a_dec_t0[19], we_a_dec_t0[19], we_a_dec_t0[19], we_a_dec_t0[19], we_a_dec_t0[19], we_a_dec_t0[19] };
  assign _0082_ = _0283_ & { we_a_dec_t0[18], we_a_dec_t0[18], we_a_dec_t0[18], we_a_dec_t0[18], we_a_dec_t0[18], we_a_dec_t0[18], we_a_dec_t0[18], we_a_dec_t0[18], we_a_dec_t0[18], we_a_dec_t0[18], we_a_dec_t0[18], we_a_dec_t0[18], we_a_dec_t0[18], we_a_dec_t0[18], we_a_dec_t0[18], we_a_dec_t0[18], we_a_dec_t0[18], we_a_dec_t0[18], we_a_dec_t0[18], we_a_dec_t0[18], we_a_dec_t0[18], we_a_dec_t0[18], we_a_dec_t0[18], we_a_dec_t0[18], we_a_dec_t0[18], we_a_dec_t0[18], we_a_dec_t0[18], we_a_dec_t0[18], we_a_dec_t0[18], we_a_dec_t0[18], we_a_dec_t0[18], we_a_dec_t0[18] };
  assign _0085_ = _0287_ & { we_a_dec_t0[17], we_a_dec_t0[17], we_a_dec_t0[17], we_a_dec_t0[17], we_a_dec_t0[17], we_a_dec_t0[17], we_a_dec_t0[17], we_a_dec_t0[17], we_a_dec_t0[17], we_a_dec_t0[17], we_a_dec_t0[17], we_a_dec_t0[17], we_a_dec_t0[17], we_a_dec_t0[17], we_a_dec_t0[17], we_a_dec_t0[17], we_a_dec_t0[17], we_a_dec_t0[17], we_a_dec_t0[17], we_a_dec_t0[17], we_a_dec_t0[17], we_a_dec_t0[17], we_a_dec_t0[17], we_a_dec_t0[17], we_a_dec_t0[17], we_a_dec_t0[17], we_a_dec_t0[17], we_a_dec_t0[17], we_a_dec_t0[17], we_a_dec_t0[17], we_a_dec_t0[17], we_a_dec_t0[17] };
  assign _0088_ = _0291_ & { we_a_dec_t0[16], we_a_dec_t0[16], we_a_dec_t0[16], we_a_dec_t0[16], we_a_dec_t0[16], we_a_dec_t0[16], we_a_dec_t0[16], we_a_dec_t0[16], we_a_dec_t0[16], we_a_dec_t0[16], we_a_dec_t0[16], we_a_dec_t0[16], we_a_dec_t0[16], we_a_dec_t0[16], we_a_dec_t0[16], we_a_dec_t0[16], we_a_dec_t0[16], we_a_dec_t0[16], we_a_dec_t0[16], we_a_dec_t0[16], we_a_dec_t0[16], we_a_dec_t0[16], we_a_dec_t0[16], we_a_dec_t0[16], we_a_dec_t0[16], we_a_dec_t0[16], we_a_dec_t0[16], we_a_dec_t0[16], we_a_dec_t0[16], we_a_dec_t0[16], we_a_dec_t0[16], we_a_dec_t0[16] };
  assign _0091_ = _0295_ & { we_a_dec_t0[15], we_a_dec_t0[15], we_a_dec_t0[15], we_a_dec_t0[15], we_a_dec_t0[15], we_a_dec_t0[15], we_a_dec_t0[15], we_a_dec_t0[15], we_a_dec_t0[15], we_a_dec_t0[15], we_a_dec_t0[15], we_a_dec_t0[15], we_a_dec_t0[15], we_a_dec_t0[15], we_a_dec_t0[15], we_a_dec_t0[15], we_a_dec_t0[15], we_a_dec_t0[15], we_a_dec_t0[15], we_a_dec_t0[15], we_a_dec_t0[15], we_a_dec_t0[15], we_a_dec_t0[15], we_a_dec_t0[15], we_a_dec_t0[15], we_a_dec_t0[15], we_a_dec_t0[15], we_a_dec_t0[15], we_a_dec_t0[15], we_a_dec_t0[15], we_a_dec_t0[15], we_a_dec_t0[15] };
  assign _0094_ = _0299_ & { we_a_dec_t0[14], we_a_dec_t0[14], we_a_dec_t0[14], we_a_dec_t0[14], we_a_dec_t0[14], we_a_dec_t0[14], we_a_dec_t0[14], we_a_dec_t0[14], we_a_dec_t0[14], we_a_dec_t0[14], we_a_dec_t0[14], we_a_dec_t0[14], we_a_dec_t0[14], we_a_dec_t0[14], we_a_dec_t0[14], we_a_dec_t0[14], we_a_dec_t0[14], we_a_dec_t0[14], we_a_dec_t0[14], we_a_dec_t0[14], we_a_dec_t0[14], we_a_dec_t0[14], we_a_dec_t0[14], we_a_dec_t0[14], we_a_dec_t0[14], we_a_dec_t0[14], we_a_dec_t0[14], we_a_dec_t0[14], we_a_dec_t0[14], we_a_dec_t0[14], we_a_dec_t0[14], we_a_dec_t0[14] };
  assign _0097_ = _0303_ & { we_a_dec_t0[13], we_a_dec_t0[13], we_a_dec_t0[13], we_a_dec_t0[13], we_a_dec_t0[13], we_a_dec_t0[13], we_a_dec_t0[13], we_a_dec_t0[13], we_a_dec_t0[13], we_a_dec_t0[13], we_a_dec_t0[13], we_a_dec_t0[13], we_a_dec_t0[13], we_a_dec_t0[13], we_a_dec_t0[13], we_a_dec_t0[13], we_a_dec_t0[13], we_a_dec_t0[13], we_a_dec_t0[13], we_a_dec_t0[13], we_a_dec_t0[13], we_a_dec_t0[13], we_a_dec_t0[13], we_a_dec_t0[13], we_a_dec_t0[13], we_a_dec_t0[13], we_a_dec_t0[13], we_a_dec_t0[13], we_a_dec_t0[13], we_a_dec_t0[13], we_a_dec_t0[13], we_a_dec_t0[13] };
  assign _0100_ = _0307_ & { we_a_dec_t0[12], we_a_dec_t0[12], we_a_dec_t0[12], we_a_dec_t0[12], we_a_dec_t0[12], we_a_dec_t0[12], we_a_dec_t0[12], we_a_dec_t0[12], we_a_dec_t0[12], we_a_dec_t0[12], we_a_dec_t0[12], we_a_dec_t0[12], we_a_dec_t0[12], we_a_dec_t0[12], we_a_dec_t0[12], we_a_dec_t0[12], we_a_dec_t0[12], we_a_dec_t0[12], we_a_dec_t0[12], we_a_dec_t0[12], we_a_dec_t0[12], we_a_dec_t0[12], we_a_dec_t0[12], we_a_dec_t0[12], we_a_dec_t0[12], we_a_dec_t0[12], we_a_dec_t0[12], we_a_dec_t0[12], we_a_dec_t0[12], we_a_dec_t0[12], we_a_dec_t0[12], we_a_dec_t0[12] };
  assign _0103_ = _0311_ & { we_a_dec_t0[11], we_a_dec_t0[11], we_a_dec_t0[11], we_a_dec_t0[11], we_a_dec_t0[11], we_a_dec_t0[11], we_a_dec_t0[11], we_a_dec_t0[11], we_a_dec_t0[11], we_a_dec_t0[11], we_a_dec_t0[11], we_a_dec_t0[11], we_a_dec_t0[11], we_a_dec_t0[11], we_a_dec_t0[11], we_a_dec_t0[11], we_a_dec_t0[11], we_a_dec_t0[11], we_a_dec_t0[11], we_a_dec_t0[11], we_a_dec_t0[11], we_a_dec_t0[11], we_a_dec_t0[11], we_a_dec_t0[11], we_a_dec_t0[11], we_a_dec_t0[11], we_a_dec_t0[11], we_a_dec_t0[11], we_a_dec_t0[11], we_a_dec_t0[11], we_a_dec_t0[11], we_a_dec_t0[11] };
  assign _0106_ = _0315_ & { we_a_dec_t0[10], we_a_dec_t0[10], we_a_dec_t0[10], we_a_dec_t0[10], we_a_dec_t0[10], we_a_dec_t0[10], we_a_dec_t0[10], we_a_dec_t0[10], we_a_dec_t0[10], we_a_dec_t0[10], we_a_dec_t0[10], we_a_dec_t0[10], we_a_dec_t0[10], we_a_dec_t0[10], we_a_dec_t0[10], we_a_dec_t0[10], we_a_dec_t0[10], we_a_dec_t0[10], we_a_dec_t0[10], we_a_dec_t0[10], we_a_dec_t0[10], we_a_dec_t0[10], we_a_dec_t0[10], we_a_dec_t0[10], we_a_dec_t0[10], we_a_dec_t0[10], we_a_dec_t0[10], we_a_dec_t0[10], we_a_dec_t0[10], we_a_dec_t0[10], we_a_dec_t0[10], we_a_dec_t0[10] };
  assign _0109_ = _0319_ & { we_a_dec_t0[9], we_a_dec_t0[9], we_a_dec_t0[9], we_a_dec_t0[9], we_a_dec_t0[9], we_a_dec_t0[9], we_a_dec_t0[9], we_a_dec_t0[9], we_a_dec_t0[9], we_a_dec_t0[9], we_a_dec_t0[9], we_a_dec_t0[9], we_a_dec_t0[9], we_a_dec_t0[9], we_a_dec_t0[9], we_a_dec_t0[9], we_a_dec_t0[9], we_a_dec_t0[9], we_a_dec_t0[9], we_a_dec_t0[9], we_a_dec_t0[9], we_a_dec_t0[9], we_a_dec_t0[9], we_a_dec_t0[9], we_a_dec_t0[9], we_a_dec_t0[9], we_a_dec_t0[9], we_a_dec_t0[9], we_a_dec_t0[9], we_a_dec_t0[9], we_a_dec_t0[9], we_a_dec_t0[9] };
  assign _0112_ = _0323_ & { we_a_dec_t0[8], we_a_dec_t0[8], we_a_dec_t0[8], we_a_dec_t0[8], we_a_dec_t0[8], we_a_dec_t0[8], we_a_dec_t0[8], we_a_dec_t0[8], we_a_dec_t0[8], we_a_dec_t0[8], we_a_dec_t0[8], we_a_dec_t0[8], we_a_dec_t0[8], we_a_dec_t0[8], we_a_dec_t0[8], we_a_dec_t0[8], we_a_dec_t0[8], we_a_dec_t0[8], we_a_dec_t0[8], we_a_dec_t0[8], we_a_dec_t0[8], we_a_dec_t0[8], we_a_dec_t0[8], we_a_dec_t0[8], we_a_dec_t0[8], we_a_dec_t0[8], we_a_dec_t0[8], we_a_dec_t0[8], we_a_dec_t0[8], we_a_dec_t0[8], we_a_dec_t0[8], we_a_dec_t0[8] };
  assign _0115_ = _0327_ & { we_a_dec_t0[7], we_a_dec_t0[7], we_a_dec_t0[7], we_a_dec_t0[7], we_a_dec_t0[7], we_a_dec_t0[7], we_a_dec_t0[7], we_a_dec_t0[7], we_a_dec_t0[7], we_a_dec_t0[7], we_a_dec_t0[7], we_a_dec_t0[7], we_a_dec_t0[7], we_a_dec_t0[7], we_a_dec_t0[7], we_a_dec_t0[7], we_a_dec_t0[7], we_a_dec_t0[7], we_a_dec_t0[7], we_a_dec_t0[7], we_a_dec_t0[7], we_a_dec_t0[7], we_a_dec_t0[7], we_a_dec_t0[7], we_a_dec_t0[7], we_a_dec_t0[7], we_a_dec_t0[7], we_a_dec_t0[7], we_a_dec_t0[7], we_a_dec_t0[7], we_a_dec_t0[7], we_a_dec_t0[7] };
  assign _0118_ = _0331_ & { we_a_dec_t0[6], we_a_dec_t0[6], we_a_dec_t0[6], we_a_dec_t0[6], we_a_dec_t0[6], we_a_dec_t0[6], we_a_dec_t0[6], we_a_dec_t0[6], we_a_dec_t0[6], we_a_dec_t0[6], we_a_dec_t0[6], we_a_dec_t0[6], we_a_dec_t0[6], we_a_dec_t0[6], we_a_dec_t0[6], we_a_dec_t0[6], we_a_dec_t0[6], we_a_dec_t0[6], we_a_dec_t0[6], we_a_dec_t0[6], we_a_dec_t0[6], we_a_dec_t0[6], we_a_dec_t0[6], we_a_dec_t0[6], we_a_dec_t0[6], we_a_dec_t0[6], we_a_dec_t0[6], we_a_dec_t0[6], we_a_dec_t0[6], we_a_dec_t0[6], we_a_dec_t0[6], we_a_dec_t0[6] };
  assign _0121_ = _0335_ & { we_a_dec_t0[5], we_a_dec_t0[5], we_a_dec_t0[5], we_a_dec_t0[5], we_a_dec_t0[5], we_a_dec_t0[5], we_a_dec_t0[5], we_a_dec_t0[5], we_a_dec_t0[5], we_a_dec_t0[5], we_a_dec_t0[5], we_a_dec_t0[5], we_a_dec_t0[5], we_a_dec_t0[5], we_a_dec_t0[5], we_a_dec_t0[5], we_a_dec_t0[5], we_a_dec_t0[5], we_a_dec_t0[5], we_a_dec_t0[5], we_a_dec_t0[5], we_a_dec_t0[5], we_a_dec_t0[5], we_a_dec_t0[5], we_a_dec_t0[5], we_a_dec_t0[5], we_a_dec_t0[5], we_a_dec_t0[5], we_a_dec_t0[5], we_a_dec_t0[5], we_a_dec_t0[5], we_a_dec_t0[5] };
  assign _0124_ = _0339_ & { we_a_dec_t0[4], we_a_dec_t0[4], we_a_dec_t0[4], we_a_dec_t0[4], we_a_dec_t0[4], we_a_dec_t0[4], we_a_dec_t0[4], we_a_dec_t0[4], we_a_dec_t0[4], we_a_dec_t0[4], we_a_dec_t0[4], we_a_dec_t0[4], we_a_dec_t0[4], we_a_dec_t0[4], we_a_dec_t0[4], we_a_dec_t0[4], we_a_dec_t0[4], we_a_dec_t0[4], we_a_dec_t0[4], we_a_dec_t0[4], we_a_dec_t0[4], we_a_dec_t0[4], we_a_dec_t0[4], we_a_dec_t0[4], we_a_dec_t0[4], we_a_dec_t0[4], we_a_dec_t0[4], we_a_dec_t0[4], we_a_dec_t0[4], we_a_dec_t0[4], we_a_dec_t0[4], we_a_dec_t0[4] };
  assign _0127_ = _0343_ & { we_a_dec_t0[3], we_a_dec_t0[3], we_a_dec_t0[3], we_a_dec_t0[3], we_a_dec_t0[3], we_a_dec_t0[3], we_a_dec_t0[3], we_a_dec_t0[3], we_a_dec_t0[3], we_a_dec_t0[3], we_a_dec_t0[3], we_a_dec_t0[3], we_a_dec_t0[3], we_a_dec_t0[3], we_a_dec_t0[3], we_a_dec_t0[3], we_a_dec_t0[3], we_a_dec_t0[3], we_a_dec_t0[3], we_a_dec_t0[3], we_a_dec_t0[3], we_a_dec_t0[3], we_a_dec_t0[3], we_a_dec_t0[3], we_a_dec_t0[3], we_a_dec_t0[3], we_a_dec_t0[3], we_a_dec_t0[3], we_a_dec_t0[3], we_a_dec_t0[3], we_a_dec_t0[3], we_a_dec_t0[3] };
  assign _0224_ = _0035_ | _0036_;
  assign _0228_ = _0038_ | _0039_;
  assign _0232_ = _0041_ | _0042_;
  assign _0236_ = _0044_ | _0045_;
  assign _0240_ = _0047_ | _0048_;
  assign _0244_ = _0050_ | _0051_;
  assign _0248_ = _0053_ | _0054_;
  assign _0252_ = _0056_ | _0057_;
  assign _0256_ = _0059_ | _0060_;
  assign _0260_ = _0062_ | _0063_;
  assign _0264_ = _0065_ | _0066_;
  assign _0268_ = _0068_ | _0069_;
  assign _0272_ = _0071_ | _0072_;
  assign _0276_ = _0074_ | _0075_;
  assign _0280_ = _0077_ | _0078_;
  assign _0284_ = _0080_ | _0081_;
  assign _0288_ = _0083_ | _0084_;
  assign _0292_ = _0086_ | _0087_;
  assign _0296_ = _0089_ | _0090_;
  assign _0300_ = _0092_ | _0093_;
  assign _0304_ = _0095_ | _0096_;
  assign _0308_ = _0098_ | _0099_;
  assign _0312_ = _0101_ | _0102_;
  assign _0316_ = _0104_ | _0105_;
  assign _0320_ = _0107_ | _0108_;
  assign _0324_ = _0110_ | _0111_;
  assign _0328_ = _0113_ | _0114_;
  assign _0332_ = _0116_ | _0117_;
  assign _0336_ = _0119_ | _0120_;
  assign _0340_ = _0122_ | _0123_;
  assign _0344_ = _0125_ | _0126_;
  assign _0225_ = _0224_ | _0037_;
  assign _0229_ = _0228_ | _0040_;
  assign _0233_ = _0232_ | _0043_;
  assign _0237_ = _0236_ | _0046_;
  assign _0241_ = _0240_ | _0049_;
  assign _0245_ = _0244_ | _0052_;
  assign _0249_ = _0248_ | _0055_;
  assign _0253_ = _0252_ | _0058_;
  assign _0257_ = _0256_ | _0061_;
  assign _0261_ = _0260_ | _0064_;
  assign _0265_ = _0264_ | _0067_;
  assign _0269_ = _0268_ | _0070_;
  assign _0273_ = _0272_ | _0073_;
  assign _0277_ = _0276_ | _0076_;
  assign _0281_ = _0280_ | _0079_;
  assign _0285_ = _0284_ | _0082_;
  assign _0289_ = _0288_ | _0085_;
  assign _0293_ = _0292_ | _0088_;
  assign _0297_ = _0296_ | _0091_;
  assign _0301_ = _0300_ | _0094_;
  assign _0305_ = _0304_ | _0097_;
  assign _0309_ = _0308_ | _0100_;
  assign _0313_ = _0312_ | _0103_;
  assign _0317_ = _0316_ | _0106_;
  assign _0321_ = _0320_ | _0109_;
  assign _0325_ = _0324_ | _0112_;
  assign _0329_ = _0328_ | _0115_;
  assign _0333_ = _0332_ | _0118_;
  assign _0337_ = _0336_ | _0121_;
  assign _0341_ = _0340_ | _0124_;
  assign _0345_ = _0344_ | _0127_;
  reg [31:0] _0782_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) _0782_ <= 32'd0;
    else _0782_ <= _0225_;
  assign rf_reg_t0[63:32] = _0782_;
  reg [31:0] _0783_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) _0783_ <= 32'd0;
    else _0783_ <= _0229_;
  assign rf_reg_t0[95:64] = _0783_;
  reg [31:0] _0784_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) _0784_ <= 32'd0;
    else _0784_ <= _0233_;
  assign rf_reg_t0[1023:992] = _0784_;
  reg [31:0] _0785_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) _0785_ <= 32'd0;
    else _0785_ <= _0237_;
  assign rf_reg_t0[991:960] = _0785_;
  reg [31:0] _0786_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) _0786_ <= 32'd0;
    else _0786_ <= _0241_;
  assign rf_reg_t0[959:928] = _0786_;
  reg [31:0] _0787_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) _0787_ <= 32'd0;
    else _0787_ <= _0245_;
  assign rf_reg_t0[927:896] = _0787_;
  reg [31:0] _0788_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) _0788_ <= 32'd0;
    else _0788_ <= _0249_;
  assign rf_reg_t0[895:864] = _0788_;
  reg [31:0] _0789_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) _0789_ <= 32'd0;
    else _0789_ <= _0253_;
  assign rf_reg_t0[863:832] = _0789_;
  reg [31:0] _0790_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) _0790_ <= 32'd0;
    else _0790_ <= _0257_;
  assign rf_reg_t0[831:800] = _0790_;
  reg [31:0] _0791_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) _0791_ <= 32'd0;
    else _0791_ <= _0261_;
  assign rf_reg_t0[799:768] = _0791_;
  reg [31:0] _0792_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) _0792_ <= 32'd0;
    else _0792_ <= _0265_;
  assign rf_reg_t0[767:736] = _0792_;
  reg [31:0] _0793_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) _0793_ <= 32'd0;
    else _0793_ <= _0269_;
  assign rf_reg_t0[735:704] = _0793_;
  reg [31:0] _0794_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) _0794_ <= 32'd0;
    else _0794_ <= _0273_;
  assign rf_reg_t0[703:672] = _0794_;
  reg [31:0] _0795_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) _0795_ <= 32'd0;
    else _0795_ <= _0277_;
  assign rf_reg_t0[671:640] = _0795_;
  reg [31:0] _0796_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) _0796_ <= 32'd0;
    else _0796_ <= _0281_;
  assign rf_reg_t0[639:608] = _0796_;
  reg [31:0] _0797_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) _0797_ <= 32'd0;
    else _0797_ <= _0285_;
  assign rf_reg_t0[607:576] = _0797_;
  reg [31:0] _0798_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) _0798_ <= 32'd0;
    else _0798_ <= _0289_;
  assign rf_reg_t0[575:544] = _0798_;
  reg [31:0] _0799_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) _0799_ <= 32'd0;
    else _0799_ <= _0293_;
  assign rf_reg_t0[543:512] = _0799_;
  reg [31:0] _0800_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) _0800_ <= 32'd0;
    else _0800_ <= _0297_;
  assign rf_reg_t0[511:480] = _0800_;
  reg [31:0] _0801_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) _0801_ <= 32'd0;
    else _0801_ <= _0301_;
  assign rf_reg_t0[479:448] = _0801_;
  reg [31:0] _0802_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) _0802_ <= 32'd0;
    else _0802_ <= _0305_;
  assign rf_reg_t0[447:416] = _0802_;
  reg [31:0] _0803_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) _0803_ <= 32'd0;
    else _0803_ <= _0309_;
  assign rf_reg_t0[415:384] = _0803_;
  reg [31:0] _0804_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) _0804_ <= 32'd0;
    else _0804_ <= _0313_;
  assign rf_reg_t0[383:352] = _0804_;
  reg [31:0] _0805_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) _0805_ <= 32'd0;
    else _0805_ <= _0317_;
  assign rf_reg_t0[351:320] = _0805_;
  reg [31:0] _0806_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) _0806_ <= 32'd0;
    else _0806_ <= _0321_;
  assign rf_reg_t0[319:288] = _0806_;
  reg [31:0] _0807_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) _0807_ <= 32'd0;
    else _0807_ <= _0325_;
  assign rf_reg_t0[287:256] = _0807_;
  reg [31:0] _0808_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) _0808_ <= 32'd0;
    else _0808_ <= _0329_;
  assign rf_reg_t0[255:224] = _0808_;
  reg [31:0] _0809_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) _0809_ <= 32'd0;
    else _0809_ <= _0333_;
  assign rf_reg_t0[223:192] = _0809_;
  reg [31:0] _0810_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) _0810_ <= 32'd0;
    else _0810_ <= _0337_;
  assign rf_reg_t0[191:160] = _0810_;
  reg [31:0] _0811_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) _0811_ <= 32'd0;
    else _0811_ <= _0341_;
  assign rf_reg_t0[159:128] = _0811_;
  reg [31:0] _0812_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) _0812_ <= 32'd0;
    else _0812_ <= _0345_;
  assign rf_reg_t0[127:96] = _0812_;
  assign _0032_ = | waddr_a_i_t0;
  assign _0031_ = ~ waddr_a_i_t0;
  assign _0128_ = waddr_a_i & _0031_;
  assign _0129_ = 5'h01 & _0031_;
  assign _0130_ = 5'h02 & _0031_;
  assign _0131_ = 5'h03 & _0031_;
  assign _0132_ = 5'h04 & _0031_;
  assign _0133_ = 5'h05 & _0031_;
  assign _0134_ = 5'h06 & _0031_;
  assign _0135_ = 5'h07 & _0031_;
  assign _0136_ = 5'h08 & _0031_;
  assign _0137_ = 5'h09 & _0031_;
  assign _0138_ = 5'h0a & _0031_;
  assign _0139_ = 5'h0b & _0031_;
  assign _0140_ = 5'h0c & _0031_;
  assign _0141_ = 5'h0d & _0031_;
  assign _0142_ = 5'h0e & _0031_;
  assign _0143_ = 5'h0f & _0031_;
  assign _0144_ = 5'h10 & _0031_;
  assign _0145_ = 5'h11 & _0031_;
  assign _0146_ = 5'h12 & _0031_;
  assign _0147_ = 5'h13 & _0031_;
  assign _0148_ = 5'h14 & _0031_;
  assign _0149_ = 5'h15 & _0031_;
  assign _0150_ = 5'h16 & _0031_;
  assign _0151_ = 5'h17 & _0031_;
  assign _0152_ = 5'h18 & _0031_;
  assign _0153_ = 5'h19 & _0031_;
  assign _0154_ = 5'h1a & _0031_;
  assign _0155_ = 5'h1b & _0031_;
  assign _0156_ = 5'h1c & _0031_;
  assign _0157_ = 5'h1d & _0031_;
  assign _0158_ = 5'h1e & _0031_;
  assign _0159_ = 5'h1f & _0031_;
  assign _0408_ = _0128_ == _0129_;
  assign _0409_ = _0128_ == _0130_;
  assign _0410_ = _0128_ == _0131_;
  assign _0411_ = _0128_ == _0132_;
  assign _0412_ = _0128_ == _0133_;
  assign _0413_ = _0128_ == _0134_;
  assign _0414_ = _0128_ == _0135_;
  assign _0415_ = _0128_ == _0136_;
  assign _0416_ = _0128_ == _0137_;
  assign _0417_ = _0128_ == _0138_;
  assign _0418_ = _0128_ == _0139_;
  assign _0419_ = _0128_ == _0140_;
  assign _0420_ = _0128_ == _0141_;
  assign _0421_ = _0128_ == _0142_;
  assign _0422_ = _0128_ == _0143_;
  assign _0423_ = _0128_ == _0144_;
  assign _0424_ = _0128_ == _0145_;
  assign _0425_ = _0128_ == _0146_;
  assign _0426_ = _0128_ == _0147_;
  assign _0427_ = _0128_ == _0148_;
  assign _0428_ = _0128_ == _0149_;
  assign _0429_ = _0128_ == _0150_;
  assign _0430_ = _0128_ == _0151_;
  assign _0431_ = _0128_ == _0152_;
  assign _0432_ = _0128_ == _0153_;
  assign _0433_ = _0128_ == _0154_;
  assign _0434_ = _0128_ == _0155_;
  assign _0435_ = _0128_ == _0156_;
  assign _0436_ = _0128_ == _0157_;
  assign _0437_ = _0128_ == _0158_;
  assign _0438_ = _0128_ == _0159_;
  assign _0442_ = _0408_ & _0032_;
  assign _0444_ = _0409_ & _0032_;
  assign _0446_ = _0410_ & _0032_;
  assign _0448_ = _0411_ & _0032_;
  assign _0450_ = _0412_ & _0032_;
  assign _0452_ = _0413_ & _0032_;
  assign _0454_ = _0414_ & _0032_;
  assign _0456_ = _0415_ & _0032_;
  assign _0458_ = _0416_ & _0032_;
  assign _0460_ = _0417_ & _0032_;
  assign _0462_ = _0418_ & _0032_;
  assign _0464_ = _0419_ & _0032_;
  assign _0466_ = _0420_ & _0032_;
  assign _0468_ = _0421_ & _0032_;
  assign _0470_ = _0422_ & _0032_;
  assign _0472_ = _0423_ & _0032_;
  assign _0474_ = _0424_ & _0032_;
  assign _0476_ = _0425_ & _0032_;
  assign _0478_ = _0426_ & _0032_;
  assign _0480_ = _0427_ & _0032_;
  assign _0482_ = _0428_ & _0032_;
  assign _0484_ = _0429_ & _0032_;
  assign _0486_ = _0430_ & _0032_;
  assign _0488_ = _0431_ & _0032_;
  assign _0490_ = _0432_ & _0032_;
  assign _0492_ = _0433_ & _0032_;
  assign _0494_ = _0434_ & _0032_;
  assign _0496_ = _0435_ & _0032_;
  assign _0498_ = _0436_ & _0032_;
  assign _0500_ = _0437_ & _0032_;
  assign _0502_ = _0438_ & _0032_;
  reg [31:0] _0909_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) _0909_ <= 32'd0;
    else if (we_a_dec[1]) _0909_ <= wdata_a_i;
  assign rf_reg[63:32] = _0909_;
  reg [31:0] _0910_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) _0910_ <= 32'd0;
    else if (we_a_dec[2]) _0910_ <= wdata_a_i;
  assign rf_reg[95:64] = _0910_;
  reg [31:0] _0911_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) _0911_ <= 32'd0;
    else if (we_a_dec[31]) _0911_ <= wdata_a_i;
  assign rf_reg[1023:992] = _0911_;
  reg [31:0] _0912_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) _0912_ <= 32'd0;
    else if (we_a_dec[30]) _0912_ <= wdata_a_i;
  assign rf_reg[991:960] = _0912_;
  reg [31:0] _0913_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) _0913_ <= 32'd0;
    else if (we_a_dec[29]) _0913_ <= wdata_a_i;
  assign rf_reg[959:928] = _0913_;
  reg [31:0] _0914_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) _0914_ <= 32'd0;
    else if (we_a_dec[28]) _0914_ <= wdata_a_i;
  assign rf_reg[927:896] = _0914_;
  reg [31:0] _0915_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) _0915_ <= 32'd0;
    else if (we_a_dec[27]) _0915_ <= wdata_a_i;
  assign rf_reg[895:864] = _0915_;
  reg [31:0] _0916_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) _0916_ <= 32'd0;
    else if (we_a_dec[26]) _0916_ <= wdata_a_i;
  assign rf_reg[863:832] = _0916_;
  reg [31:0] _0917_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) _0917_ <= 32'd0;
    else if (we_a_dec[25]) _0917_ <= wdata_a_i;
  assign rf_reg[831:800] = _0917_;
  reg [31:0] _0918_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) _0918_ <= 32'd0;
    else if (we_a_dec[24]) _0918_ <= wdata_a_i;
  assign rf_reg[799:768] = _0918_;
  reg [31:0] _0919_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) _0919_ <= 32'd0;
    else if (we_a_dec[23]) _0919_ <= wdata_a_i;
  assign rf_reg[767:736] = _0919_;
  reg [31:0] _0920_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) _0920_ <= 32'd0;
    else if (we_a_dec[22]) _0920_ <= wdata_a_i;
  assign rf_reg[735:704] = _0920_;
  reg [31:0] _0921_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) _0921_ <= 32'd0;
    else if (we_a_dec[21]) _0921_ <= wdata_a_i;
  assign rf_reg[703:672] = _0921_;
  reg [31:0] _0922_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) _0922_ <= 32'd0;
    else if (we_a_dec[20]) _0922_ <= wdata_a_i;
  assign rf_reg[671:640] = _0922_;
  reg [31:0] _0923_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) _0923_ <= 32'd0;
    else if (we_a_dec[19]) _0923_ <= wdata_a_i;
  assign rf_reg[639:608] = _0923_;
  reg [31:0] _0924_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) _0924_ <= 32'd0;
    else if (we_a_dec[18]) _0924_ <= wdata_a_i;
  assign rf_reg[607:576] = _0924_;
  reg [31:0] _0925_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) _0925_ <= 32'd0;
    else if (we_a_dec[17]) _0925_ <= wdata_a_i;
  assign rf_reg[575:544] = _0925_;
  reg [31:0] _0926_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) _0926_ <= 32'd0;
    else if (we_a_dec[16]) _0926_ <= wdata_a_i;
  assign rf_reg[543:512] = _0926_;
  reg [31:0] _0927_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) _0927_ <= 32'd0;
    else if (we_a_dec[15]) _0927_ <= wdata_a_i;
  assign rf_reg[511:480] = _0927_;
  reg [31:0] _0928_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) _0928_ <= 32'd0;
    else if (we_a_dec[14]) _0928_ <= wdata_a_i;
  assign rf_reg[479:448] = _0928_;
  reg [31:0] _0929_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) _0929_ <= 32'd0;
    else if (we_a_dec[13]) _0929_ <= wdata_a_i;
  assign rf_reg[447:416] = _0929_;
  reg [31:0] _0930_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) _0930_ <= 32'd0;
    else if (we_a_dec[12]) _0930_ <= wdata_a_i;
  assign rf_reg[415:384] = _0930_;
  reg [31:0] _0931_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) _0931_ <= 32'd0;
    else if (we_a_dec[11]) _0931_ <= wdata_a_i;
  assign rf_reg[383:352] = _0931_;
  reg [31:0] _0932_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) _0932_ <= 32'd0;
    else if (we_a_dec[10]) _0932_ <= wdata_a_i;
  assign rf_reg[351:320] = _0932_;
  reg [31:0] _0933_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) _0933_ <= 32'd0;
    else if (we_a_dec[9]) _0933_ <= wdata_a_i;
  assign rf_reg[319:288] = _0933_;
  reg [31:0] _0934_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) _0934_ <= 32'd0;
    else if (we_a_dec[8]) _0934_ <= wdata_a_i;
  assign rf_reg[287:256] = _0934_;
  reg [31:0] _0935_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) _0935_ <= 32'd0;
    else if (we_a_dec[7]) _0935_ <= wdata_a_i;
  assign rf_reg[255:224] = _0935_;
  reg [31:0] _0936_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) _0936_ <= 32'd0;
    else if (we_a_dec[6]) _0936_ <= wdata_a_i;
  assign rf_reg[223:192] = _0936_;
  reg [31:0] _0937_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) _0937_ <= 32'd0;
    else if (we_a_dec[5]) _0937_ <= wdata_a_i;
  assign rf_reg[191:160] = _0937_;
  reg [31:0] _0938_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) _0938_ <= 32'd0;
    else if (we_a_dec[4]) _0938_ <= wdata_a_i;
  assign rf_reg[159:128] = _0938_;
  reg [31:0] _0939_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) _0939_ <= 32'd0;
    else if (we_a_dec[3]) _0939_ <= wdata_a_i;
  assign rf_reg[127:96] = _0939_;
  assign _0346_ = _0442_ | _0441_;
  assign _0347_ = _0444_ | _0443_;
  assign _0348_ = _0446_ | _0445_;
  assign _0349_ = _0448_ | _0447_;
  assign _0350_ = _0450_ | _0449_;
  assign _0351_ = _0452_ | _0451_;
  assign _0352_ = _0454_ | _0453_;
  assign _0353_ = _0456_ | _0455_;
  assign _0354_ = _0458_ | _0457_;
  assign _0355_ = _0460_ | _0459_;
  assign _0356_ = _0462_ | _0461_;
  assign _0357_ = _0464_ | _0463_;
  assign _0358_ = _0466_ | _0465_;
  assign _0359_ = _0468_ | _0467_;
  assign _0360_ = _0470_ | _0469_;
  assign _0361_ = _0472_ | _0471_;
  assign _0362_ = _0474_ | _0473_;
  assign _0363_ = _0476_ | _0475_;
  assign _0364_ = _0478_ | _0477_;
  assign _0365_ = _0480_ | _0479_;
  assign _0366_ = _0482_ | _0481_;
  assign _0367_ = _0484_ | _0483_;
  assign _0368_ = _0486_ | _0485_;
  assign _0369_ = _0488_ | _0487_;
  assign _0370_ = _0490_ | _0489_;
  assign _0371_ = _0492_ | _0491_;
  assign _0372_ = _0494_ | _0493_;
  assign _0373_ = _0496_ | _0495_;
  assign _0374_ = _0498_ | _0497_;
  assign _0375_ = _0500_ | _0499_;
  assign _0376_ = _0502_ | _0501_;
  assign _0160_ = we_a_i_t0 & _0346_;
  assign _0162_ = we_a_i_t0 & _0347_;
  assign _0164_ = we_a_i_t0 & _0348_;
  assign _0166_ = we_a_i_t0 & _0349_;
  assign _0168_ = we_a_i_t0 & _0350_;
  assign _0170_ = we_a_i_t0 & _0351_;
  assign _0172_ = we_a_i_t0 & _0352_;
  assign _0174_ = we_a_i_t0 & _0353_;
  assign _0176_ = we_a_i_t0 & _0354_;
  assign _0178_ = we_a_i_t0 & _0355_;
  assign _0180_ = we_a_i_t0 & _0356_;
  assign _0182_ = we_a_i_t0 & _0357_;
  assign _0184_ = we_a_i_t0 & _0358_;
  assign _0186_ = we_a_i_t0 & _0359_;
  assign _0188_ = we_a_i_t0 & _0360_;
  assign _0190_ = we_a_i_t0 & _0361_;
  assign _0192_ = we_a_i_t0 & _0362_;
  assign _0194_ = we_a_i_t0 & _0363_;
  assign _0196_ = we_a_i_t0 & _0364_;
  assign _0198_ = we_a_i_t0 & _0365_;
  assign _0200_ = we_a_i_t0 & _0366_;
  assign _0202_ = we_a_i_t0 & _0367_;
  assign _0204_ = we_a_i_t0 & _0368_;
  assign _0206_ = we_a_i_t0 & _0369_;
  assign _0208_ = we_a_i_t0 & _0370_;
  assign _0210_ = we_a_i_t0 & _0371_;
  assign _0212_ = we_a_i_t0 & _0372_;
  assign _0214_ = we_a_i_t0 & _0373_;
  assign _0216_ = we_a_i_t0 & _0374_;
  assign _0218_ = we_a_i_t0 & _0375_;
  assign _0220_ = we_a_i_t0 & _0376_;
  assign _0161_ = _0442_ & we_a_i;
  assign _0163_ = _0444_ & we_a_i;
  assign _0165_ = _0446_ & we_a_i;
  assign _0167_ = _0448_ & we_a_i;
  assign _0169_ = _0450_ & we_a_i;
  assign _0171_ = _0452_ & we_a_i;
  assign _0173_ = _0454_ & we_a_i;
  assign _0175_ = _0456_ & we_a_i;
  assign _0177_ = _0458_ & we_a_i;
  assign _0179_ = _0460_ & we_a_i;
  assign _0181_ = _0462_ & we_a_i;
  assign _0183_ = _0464_ & we_a_i;
  assign _0185_ = _0466_ & we_a_i;
  assign _0187_ = _0468_ & we_a_i;
  assign _0189_ = _0470_ & we_a_i;
  assign _0191_ = _0472_ & we_a_i;
  assign _0193_ = _0474_ & we_a_i;
  assign _0195_ = _0476_ & we_a_i;
  assign _0197_ = _0478_ & we_a_i;
  assign _0199_ = _0480_ & we_a_i;
  assign _0201_ = _0482_ & we_a_i;
  assign _0203_ = _0484_ & we_a_i;
  assign _0205_ = _0486_ & we_a_i;
  assign _0207_ = _0488_ & we_a_i;
  assign _0209_ = _0490_ & we_a_i;
  assign _0211_ = _0492_ & we_a_i;
  assign _0213_ = _0494_ & we_a_i;
  assign _0215_ = _0496_ & we_a_i;
  assign _0217_ = _0498_ & we_a_i;
  assign _0219_ = _0500_ & we_a_i;
  assign _0221_ = _0502_ & we_a_i;
  assign we_a_dec_t0[1] = _0161_ | _0160_;
  assign we_a_dec_t0[2] = _0163_ | _0162_;
  assign we_a_dec_t0[3] = _0165_ | _0164_;
  assign we_a_dec_t0[4] = _0167_ | _0166_;
  assign we_a_dec_t0[5] = _0169_ | _0168_;
  assign we_a_dec_t0[6] = _0171_ | _0170_;
  assign we_a_dec_t0[7] = _0173_ | _0172_;
  assign we_a_dec_t0[8] = _0175_ | _0174_;
  assign we_a_dec_t0[9] = _0177_ | _0176_;
  assign we_a_dec_t0[10] = _0179_ | _0178_;
  assign we_a_dec_t0[11] = _0181_ | _0180_;
  assign we_a_dec_t0[12] = _0183_ | _0182_;
  assign we_a_dec_t0[13] = _0185_ | _0184_;
  assign we_a_dec_t0[14] = _0187_ | _0186_;
  assign we_a_dec_t0[15] = _0189_ | _0188_;
  assign we_a_dec_t0[16] = _0191_ | _0190_;
  assign we_a_dec_t0[17] = _0193_ | _0192_;
  assign we_a_dec_t0[18] = _0195_ | _0194_;
  assign we_a_dec_t0[19] = _0197_ | _0196_;
  assign we_a_dec_t0[20] = _0199_ | _0198_;
  assign we_a_dec_t0[21] = _0201_ | _0200_;
  assign we_a_dec_t0[22] = _0203_ | _0202_;
  assign we_a_dec_t0[23] = _0205_ | _0204_;
  assign we_a_dec_t0[24] = _0207_ | _0206_;
  assign we_a_dec_t0[25] = _0209_ | _0208_;
  assign we_a_dec_t0[26] = _0211_ | _0210_;
  assign we_a_dec_t0[27] = _0213_ | _0212_;
  assign we_a_dec_t0[28] = _0215_ | _0214_;
  assign we_a_dec_t0[29] = _0217_ | _0216_;
  assign we_a_dec_t0[30] = _0219_ | _0218_;
  assign we_a_dec_t0[31] = _0221_ | _0220_;
  assign _0033_ = | raddr_a_i_t0;
  assign _0034_ = | raddr_b_i_t0;
  wire [1023:0] _1134_ = { rf_reg_t0[1023:32], 32'h00000000 };
  assign _0439_ = _1134_[$signed({ 22'h000000, raddr_a_i, 5'h00 }) +: 32];
  wire [1023:0] _1135_ = { rf_reg_t0[1023:32], 32'h00000000 };
  assign _0440_ = _1135_[$signed({ 22'h000000, raddr_b_i, 5'h00 }) +: 32];
  assign rdata_a_o_t0 = { _0033_, _0033_, _0033_, _0033_, _0033_, _0033_, _0033_, _0033_, _0033_, _0033_, _0033_, _0033_, _0033_, _0033_, _0033_, _0033_, _0033_, _0033_, _0033_, _0033_, _0033_, _0033_, _0033_, _0033_, _0033_, _0033_, _0033_, _0033_, _0033_, _0033_, _0033_, _0033_ } | _0439_;
  assign rdata_b_o_t0 = { _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_ } | _0440_;
  assign _0441_ = waddr_a_i == 5'h01;
  assign _0443_ = waddr_a_i == 5'h02;
  assign _0445_ = waddr_a_i == 5'h03;
  assign _0447_ = waddr_a_i == 5'h04;
  assign _0449_ = waddr_a_i == 5'h05;
  assign _0451_ = waddr_a_i == 5'h06;
  assign _0453_ = waddr_a_i == 5'h07;
  assign _0455_ = waddr_a_i == 5'h08;
  assign _0457_ = waddr_a_i == 5'h09;
  assign _0459_ = waddr_a_i == 5'h0a;
  assign _0461_ = waddr_a_i == 5'h0b;
  assign _0463_ = waddr_a_i == 5'h0c;
  assign _0465_ = waddr_a_i == 5'h0d;
  assign _0467_ = waddr_a_i == 5'h0e;
  assign _0469_ = waddr_a_i == 5'h0f;
  assign _0471_ = waddr_a_i == 5'h10;
  assign _0473_ = waddr_a_i == 5'h11;
  assign _0475_ = waddr_a_i == 5'h12;
  assign _0477_ = waddr_a_i == 5'h13;
  assign _0479_ = waddr_a_i == 5'h14;
  assign _0481_ = waddr_a_i == 5'h15;
  assign _0483_ = waddr_a_i == 5'h16;
  assign _0485_ = waddr_a_i == 5'h17;
  assign _0487_ = waddr_a_i == 5'h18;
  assign _0489_ = waddr_a_i == 5'h19;
  assign _0491_ = waddr_a_i == 5'h1a;
  assign _0493_ = waddr_a_i == 5'h1b;
  assign _0495_ = waddr_a_i == 5'h1c;
  assign _0497_ = waddr_a_i == 5'h1d;
  assign _0499_ = waddr_a_i == 5'h1e;
  assign _0501_ = waddr_a_i == 5'h1f;
  wire [1023:0] _1136_ = { rf_reg[1023:32], 32'h00000000 };
  assign rdata_a_o = _1136_[$signed({ 22'h000000, raddr_a_i, 5'h00 }) +: 32];
  wire [1023:0] _1137_ = { rf_reg[1023:32], 32'h00000000 };
  assign rdata_b_o = _1137_[$signed({ 22'h000000, raddr_b_i, 5'h00 }) +: 32];
  assign we_a_dec[1] = _0441_ ? we_a_i : 1'h0;
  assign we_a_dec[2] = _0443_ ? we_a_i : 1'h0;
  assign we_a_dec[3] = _0445_ ? we_a_i : 1'h0;
  assign we_a_dec[4] = _0447_ ? we_a_i : 1'h0;
  assign we_a_dec[5] = _0449_ ? we_a_i : 1'h0;
  assign we_a_dec[6] = _0451_ ? we_a_i : 1'h0;
  assign we_a_dec[7] = _0453_ ? we_a_i : 1'h0;
  assign we_a_dec[8] = _0455_ ? we_a_i : 1'h0;
  assign we_a_dec[9] = _0457_ ? we_a_i : 1'h0;
  assign we_a_dec[10] = _0459_ ? we_a_i : 1'h0;
  assign we_a_dec[11] = _0461_ ? we_a_i : 1'h0;
  assign we_a_dec[12] = _0463_ ? we_a_i : 1'h0;
  assign we_a_dec[13] = _0465_ ? we_a_i : 1'h0;
  assign we_a_dec[14] = _0467_ ? we_a_i : 1'h0;
  assign we_a_dec[15] = _0469_ ? we_a_i : 1'h0;
  assign we_a_dec[16] = _0471_ ? we_a_i : 1'h0;
  assign we_a_dec[17] = _0473_ ? we_a_i : 1'h0;
  assign we_a_dec[18] = _0475_ ? we_a_i : 1'h0;
  assign we_a_dec[19] = _0477_ ? we_a_i : 1'h0;
  assign we_a_dec[20] = _0479_ ? we_a_i : 1'h0;
  assign we_a_dec[21] = _0481_ ? we_a_i : 1'h0;
  assign we_a_dec[22] = _0483_ ? we_a_i : 1'h0;
  assign we_a_dec[23] = _0485_ ? we_a_i : 1'h0;
  assign we_a_dec[24] = _0487_ ? we_a_i : 1'h0;
  assign we_a_dec[25] = _0489_ ? we_a_i : 1'h0;
  assign we_a_dec[26] = _0491_ ? we_a_i : 1'h0;
  assign we_a_dec[27] = _0493_ ? we_a_i : 1'h0;
  assign we_a_dec[28] = _0495_ ? we_a_i : 1'h0;
  assign we_a_dec[29] = _0497_ ? we_a_i : 1'h0;
  assign we_a_dec[30] = _0499_ ? we_a_i : 1'h0;
  assign we_a_dec[31] = _0501_ ? we_a_i : 1'h0;
  assign rf_reg[31:0] = 32'd0;
  assign rf_reg_t0[31:0] = 32'd0;
endmodule

module paramod228b056930db4609081e7d118c0624e476409ccbauxy_ibex_if_stage (clk_i, rst_ni, boot_addr_i, req_i, instr_req_o, instr_addr_o, instr_gnt_i, instr_rvalid_i, instr_rdata_i, instr_err_i, instr_pmp_err_i, ic_tag_req_o, ic_tag_write_o, ic_tag_addr_o, ic_tag_wdata_o, ic_tag_rdata_i, ic_data_req_o, ic_data_write_o, ic_data_addr_o, ic_data_wdata_o, ic_data_rdata_i
, instr_valid_id_o, instr_new_id_o, instr_rdata_id_o, instr_rdata_alu_id_o, instr_rdata_c_id_o, instr_is_compressed_id_o, instr_bp_taken_o, instr_fetch_err_o, instr_fetch_err_plus2_o, illegal_c_insn_id_o, dummy_instr_id_o, pc_if_o, pc_id_o, instr_valid_clear_i, pc_set_i, pc_set_spec_i, pc_mux_i, nt_branch_mispredict_i, exc_pc_mux_i, exc_cause, dummy_instr_en_i
, dummy_instr_mask_i, dummy_instr_seed_en_i, dummy_instr_seed_i, icache_enable_i, icache_inval_i, branch_target_ex_i, csr_mepc_i, csr_depc_i, csr_mtvec_i, csr_mtvec_init_o, id_in_ready_i, pc_mismatch_alert_o, if_busy_o, if_busy_o_t0, id_in_ready_i_t0, icache_inval_i_t0, icache_enable_i_t0, ic_tag_write_o_t0, ic_tag_wdata_o_t0, ic_tag_req_o_t0, ic_tag_rdata_i_t0
, ic_tag_addr_o_t0, ic_data_write_o_t0, ic_data_wdata_o_t0, ic_data_req_o_t0, ic_data_rdata_i_t0, ic_data_addr_o_t0, exc_pc_mux_i_t0, exc_cause_t0, dummy_instr_seed_en_i_t0, dummy_instr_en_i_t0, csr_mtvec_init_o_t0, boot_addr_i_t0, pc_set_spec_i_t0, pc_set_i_t0, pc_mux_i_t0, pc_mismatch_alert_o_t0, pc_if_o_t0, pc_id_o_t0, nt_branch_mispredict_i_t0, instr_valid_id_o_t0, instr_valid_clear_i_t0
, instr_rdata_id_o_t0, instr_rdata_c_id_o_t0, instr_rdata_alu_id_o_t0, instr_new_id_o_t0, instr_is_compressed_id_o_t0, instr_fetch_err_plus2_o_t0, instr_fetch_err_o_t0, instr_bp_taken_o_t0, illegal_c_insn_id_o_t0, dummy_instr_seed_i_t0, dummy_instr_mask_i_t0, dummy_instr_id_o_t0, csr_mtvec_i_t0, csr_mepc_i_t0, csr_depc_i_t0, branch_target_ex_i_t0, req_i_t0, instr_rvalid_i_t0, instr_req_o_t0, instr_rdata_i_t0, instr_pmp_err_i_t0
, instr_gnt_i_t0, instr_err_i_t0, instr_addr_o_t0);
  wire signal000;
  wire signal001;
  wire signal002;
  wire signal003;
  wire signal004;
  wire signal005;
  wire signal006;
  wire signal007;
  wire signal008;
  wire signal009;
  wire signal010;
  wire [31:0] signal011;
  wire [31:0] signal012;
  wire [31:0] signal013;
  wire [31:0] signal014;
  wire [31:0] signal015;
  wire [31:0] signal016;
  wire [31:0] signal017;
  wire [2:0] signal018;
  wire signal019;
  wire signal020;
  wire [1:0] signal021;
  wire signal022;
  wire signal023;
  wire signal024;
  wire signal025;
  wire signal026;
  wire signal027;
  wire signal028;
  wire signal029;
  wire signal030;
  wire signal031;
  wire signal032;
  wire signal033;
  wire signal034;
  wire signal035;
  wire signal036;
  wire signal037;
  wire signal038;
  wire signal039;
  wire [31:0] signal040;
  wire [31:0] signal041;
  wire [31:0] signal042;
  wire signal043;
  wire signal044;
  wire signal045;
  wire signal046;
  wire signal047;
  wire signal048;
  wire [15:0] signal049;
  wire [15:0] signal050;
  wire [15:0] signal051;
  wire signal052;
  wire signal053;
  wire signal054;
  wire signal055;
  wire signal056;
  wire signal057;
  wire [31:0] signal058;
  wire [31:0] signal059;
  wire [31:0] signal060;
  wire signal061;
  wire signal062;
  wire signal063;
  wire signal064;
  wire signal065;
  wire signal066;
  wire [31:0] signal067;
  wire [31:0] signal068;
  wire [31:0] signal069;
  wire [31:0] signal070;
  wire [31:0] signal071;
  wire [31:0] signal072;
  wire [31:0] signal073;
  wire [31:0] signal074;
  wire [31:0] signal075;
  wire [31:0] signal076;
  wire [31:0] signal077;
  wire [31:0] signal078;
  wire [31:0] signal079;
  wire [31:0] signal080;
  wire [31:0] signal081;
  wire [31:0] signal082;
  wire [31:0] signal083;
  wire [31:0] signal084;
  wire [31:0] signal085;
  wire [31:0] signal086;
  wire [31:0] signal087;
  wire [2:0] signal088;
  wire signal089;
  wire signal090;
  wire signal091;
  wire [2:0] signal092;
  wire [2:0] signal093;
  wire [2:0] signal094;
  wire [2:0] signal095;
  wire [1:0] signal096;
  wire [1:0] signal097;
  wire [1:0] signal098;
  wire [1:0] signal099;
  wire signal100;
  wire signal101;
  wire signal102;
  wire signal103;
  wire signal104;
  wire signal105;
  wire signal106;
  wire signal107;
  wire signal108;
  wire [31:0] signal109;
  wire [31:0] signal110;
  wire [31:0] signal111;
  wire [31:0] signal112;
  wire signal113;
  wire signal114;
  wire signal115;
  wire signal116;
  wire signal117;
  wire signal118;
  wire signal119;
  wire signal120;
  wire [15:0] signal121;
  wire [15:0] signal122;
  wire [15:0] signal123;
  wire [15:0] signal124;
  wire signal125;
  wire signal126;
  wire signal127;
  wire signal128;
  wire signal129;
  wire signal130;
  wire signal131;
  wire signal132;
  wire [31:0] signal133;
  wire [31:0] signal134;
  wire [31:0] signal135;
  wire [31:0] signal136;
  wire signal137;
  wire signal138;
  wire [31:0] signal139;
  wire [31:0] signal140;
  wire [31:0] signal141;
  wire [31:0] signal142;
  wire [31:0] signal143;
  wire [31:0] signal144;
  wire [31:0] signal145;
  wire [31:0] signal146;
  wire [31:0] signal147;
  wire [31:0] signal148;
  wire [31:0] signal149;
  wire [31:0] signal150;
  wire [31:0] signal151;
  wire [31:0] signal152;
  wire [31:0] signal153;
  wire [31:0] signal154;
  wire [31:0] signal155;
  wire [31:0] signal156;
  wire [31:0] signal157;
  wire [31:0] signal158;
  wire [31:0] signal159;
  wire signal160;
  wire [31:0] signal161;
  wire signal162;
  wire signal163;
  wire [15:0] signal164;
  wire signal165;
  wire signal166;
  wire [31:0] signal167;
  wire [31:0] signal168;
  wire [31:0] signal169;
  wire [31:0] signal170;
  wire [31:0] signal171;
  wire [31:0] signal172;
  wire [31:0] signal173;
  wire signal174;
  wire signal175;
  wire signal176;
  wire signal177;
  wire signal178;
  wire signal179;
  wire signal180;
  wire [31:0] signal181;
  wire [31:0] signal182;
  wire [31:0] signal183;
  wire [31:0] signal184;
  wire [31:0] signal185;
  wire [31:0] signal186;
  wire [31:0] signal187;
  wire [31:0] signal188;
  wire [31:0] signal189;
  wire [31:0] signal190;
  wire signal191;
  wire signal192;
  wire signal193;
  wire signal194;
  wire signal195;
  wire signal196;
  wire signal197;
  wire signal198;
  wire signal199;
  wire signal200;
  wire signal201;
  wire signal202;
  wire signal203;
  wire signal204;
  wire signal205;
  wire signal206;
  wire signal207;
  wire signal208;
  wire signal209;
  input [31:0] boot_addr_i;
  wire [31:0] boot_addr_i;
  input [31:0] boot_addr_i_t0;
  wire [31:0] boot_addr_i_t0;
  input [31:0] branch_target_ex_i;
  wire [31:0] branch_target_ex_i;
  input [31:0] branch_target_ex_i_t0;
  wire [31:0] branch_target_ex_i_t0;
  input clk_i;
  wire clk_i;
  input [31:0] csr_depc_i;
  wire [31:0] csr_depc_i;
  input [31:0] csr_depc_i_t0;
  wire [31:0] csr_depc_i_t0;
  input [31:0] csr_mepc_i;
  wire [31:0] csr_mepc_i;
  input [31:0] csr_mepc_i_t0;
  wire [31:0] csr_mepc_i_t0;
  input [31:0] csr_mtvec_i;
  wire [31:0] csr_mtvec_i;
  input [31:0] csr_mtvec_i_t0;
  wire [31:0] csr_mtvec_i_t0;
  output csr_mtvec_init_o;
  wire csr_mtvec_init_o;
  output csr_mtvec_init_o_t0;
  wire csr_mtvec_init_o_t0;
  input dummy_instr_en_i;
  wire dummy_instr_en_i;
  input dummy_instr_en_i_t0;
  wire dummy_instr_en_i_t0;
  output dummy_instr_id_o;
  wire dummy_instr_id_o;
  output dummy_instr_id_o_t0;
  wire dummy_instr_id_o_t0;
  input [2:0] dummy_instr_mask_i;
  wire [2:0] dummy_instr_mask_i;
  input [2:0] dummy_instr_mask_i_t0;
  wire [2:0] dummy_instr_mask_i_t0;
  input dummy_instr_seed_en_i;
  wire dummy_instr_seed_en_i;
  input dummy_instr_seed_en_i_t0;
  wire dummy_instr_seed_en_i_t0;
  input [31:0] dummy_instr_seed_i;
  wire [31:0] dummy_instr_seed_i;
  input [31:0] dummy_instr_seed_i_t0;
  wire [31:0] dummy_instr_seed_i_t0;
  input [5:0] exc_cause;
  wire [5:0] exc_cause;
  input [5:0] exc_cause_t0;
  wire [5:0] exc_cause_t0;
  wire [31:0] exc_pc;
  input [1:0] exc_pc_mux_i;
  wire [1:0] exc_pc_mux_i;
  input [1:0] exc_pc_mux_i_t0;
  wire [1:0] exc_pc_mux_i_t0;
  wire [31:0] exc_pc_t0;
  wire [31:0] fetch_addr_n;
  wire [31:0] fetch_addr_n_t0;
  wire fetch_err;
  wire fetch_err_plus2;
  wire fetch_err_plus2_t0;
  wire fetch_err_t0;
  wire [31:0] fetch_rdata;
  wire [31:0] fetch_rdata_t0;
  wire fetch_valid;
  wire fetch_valid_t0;
  output [7:0] ic_data_addr_o;
  wire [7:0] ic_data_addr_o;
  output [7:0] ic_data_addr_o_t0;
  wire [7:0] ic_data_addr_o_t0;
  input [127:0] ic_data_rdata_i;
  wire [127:0] ic_data_rdata_i;
  input [127:0] ic_data_rdata_i_t0;
  wire [127:0] ic_data_rdata_i_t0;
  output [1:0] ic_data_req_o;
  wire [1:0] ic_data_req_o;
  output [1:0] ic_data_req_o_t0;
  wire [1:0] ic_data_req_o_t0;
  output [63:0] ic_data_wdata_o;
  wire [63:0] ic_data_wdata_o;
  output [63:0] ic_data_wdata_o_t0;
  wire [63:0] ic_data_wdata_o_t0;
  output ic_data_write_o;
  wire ic_data_write_o;
  output ic_data_write_o_t0;
  wire ic_data_write_o_t0;
  output [7:0] ic_tag_addr_o;
  wire [7:0] ic_tag_addr_o;
  output [7:0] ic_tag_addr_o_t0;
  wire [7:0] ic_tag_addr_o_t0;
  input [43:0] ic_tag_rdata_i;
  wire [43:0] ic_tag_rdata_i;
  input [43:0] ic_tag_rdata_i_t0;
  wire [43:0] ic_tag_rdata_i_t0;
  output [1:0] ic_tag_req_o;
  wire [1:0] ic_tag_req_o;
  output [1:0] ic_tag_req_o_t0;
  wire [1:0] ic_tag_req_o_t0;
  output [21:0] ic_tag_wdata_o;
  wire [21:0] ic_tag_wdata_o;
  output [21:0] ic_tag_wdata_o_t0;
  wire [21:0] ic_tag_wdata_o_t0;
  output ic_tag_write_o;
  wire ic_tag_write_o;
  output ic_tag_write_o_t0;
  wire ic_tag_write_o_t0;
  input icache_enable_i;
  wire icache_enable_i;
  input icache_enable_i_t0;
  wire icache_enable_i_t0;
  input icache_inval_i;
  wire icache_inval_i;
  input icache_inval_i_t0;
  wire icache_inval_i_t0;
  input id_in_ready_i;
  wire id_in_ready_i;
  input id_in_ready_i_t0;
  wire id_in_ready_i_t0;
  output if_busy_o;
  wire if_busy_o;
  output if_busy_o_t0;
  wire if_busy_o_t0;
  wire if_id_pipe_reg_we;
  wire if_id_pipe_reg_we_t0;
  wire illegal_c_insn;
  output illegal_c_insn_id_o;
  reg illegal_c_insn_id_o;
  output illegal_c_insn_id_o_t0;
  reg illegal_c_insn_id_o_t0;
  wire illegal_c_insn_t0;
  output [31:0] instr_addr_o;
  wire [31:0] instr_addr_o;
  output [31:0] instr_addr_o_t0;
  wire [31:0] instr_addr_o_t0;
  output instr_bp_taken_o;
  wire instr_bp_taken_o;
  output instr_bp_taken_o_t0;
  wire instr_bp_taken_o_t0;
  wire [31:0] instr_decompressed;
  wire [31:0] instr_decompressed_t0;
  input instr_err_i;
  wire instr_err_i;
  input instr_err_i_t0;
  wire instr_err_i_t0;
  output instr_fetch_err_o;
  reg instr_fetch_err_o;
  output instr_fetch_err_o_t0;
  reg instr_fetch_err_o_t0;
  output instr_fetch_err_plus2_o;
  reg instr_fetch_err_plus2_o;
  output instr_fetch_err_plus2_o_t0;
  reg instr_fetch_err_plus2_o_t0;
  input instr_gnt_i;
  wire instr_gnt_i;
  input instr_gnt_i_t0;
  wire instr_gnt_i_t0;
  wire instr_is_compressed;
  output instr_is_compressed_id_o;
  reg instr_is_compressed_id_o;
  output instr_is_compressed_id_o_t0;
  reg instr_is_compressed_id_o_t0;
  wire instr_is_compressed_t0;
  output instr_new_id_o;
  reg instr_new_id_o;
  output instr_new_id_o_t0;
  reg instr_new_id_o_t0;
  input instr_pmp_err_i;
  wire instr_pmp_err_i;
  input instr_pmp_err_i_t0;
  wire instr_pmp_err_i_t0;
  output [31:0] instr_rdata_alu_id_o;
  reg [31:0] instr_rdata_alu_id_o;
  output [31:0] instr_rdata_alu_id_o_t0;
  reg [31:0] instr_rdata_alu_id_o_t0;
  output [15:0] instr_rdata_c_id_o;
  reg [15:0] instr_rdata_c_id_o;
  output [15:0] instr_rdata_c_id_o_t0;
  reg [15:0] instr_rdata_c_id_o_t0;
  input [31:0] instr_rdata_i;
  wire [31:0] instr_rdata_i;
  input [31:0] instr_rdata_i_t0;
  wire [31:0] instr_rdata_i_t0;
  output [31:0] instr_rdata_id_o;
  wire [31:0] instr_rdata_id_o;
  output [31:0] instr_rdata_id_o_t0;
  wire [31:0] instr_rdata_id_o_t0;
  output instr_req_o;
  wire instr_req_o;
  output instr_req_o_t0;
  wire instr_req_o_t0;
  input instr_rvalid_i;
  wire instr_rvalid_i;
  input instr_rvalid_i_t0;
  wire instr_rvalid_i_t0;
  input instr_valid_clear_i;
  wire instr_valid_clear_i;
  input instr_valid_clear_i_t0;
  wire instr_valid_clear_i_t0;
  wire instr_valid_id_d;
  wire instr_valid_id_d_t0;
  output instr_valid_id_o;
  reg instr_valid_id_o;
  output instr_valid_id_o_t0;
  reg instr_valid_id_o_t0;
  input nt_branch_mispredict_i;
  wire nt_branch_mispredict_i;
  input nt_branch_mispredict_i_t0;
  wire nt_branch_mispredict_i_t0;
  output [31:0] pc_id_o;
  reg [31:0] pc_id_o;
  output [31:0] pc_id_o_t0;
  reg [31:0] pc_id_o_t0;
  output [31:0] pc_if_o;
  wire [31:0] pc_if_o;
  output [31:0] pc_if_o_t0;
  wire [31:0] pc_if_o_t0;
  output pc_mismatch_alert_o;
  wire pc_mismatch_alert_o;
  output pc_mismatch_alert_o_t0;
  wire pc_mismatch_alert_o_t0;
  input [2:0] pc_mux_i;
  wire [2:0] pc_mux_i;
  input [2:0] pc_mux_i_t0;
  wire [2:0] pc_mux_i_t0;
  input pc_set_i;
  wire pc_set_i;
  input pc_set_i_t0;
  wire pc_set_i_t0;
  input pc_set_spec_i;
  wire pc_set_spec_i;
  input pc_set_spec_i_t0;
  wire pc_set_spec_i_t0;
  input req_i;
  wire req_i;
  input req_i_t0;
  wire req_i_t0;
  input rst_ni;
  wire rst_ni;
  assign csr_mtvec_init_o = signal191 & pc_set_i;
  assign signal000 = fetch_valid & signal193;
  assign signal002 = if_id_pipe_reg_we & signal194;
  assign signal004 = instr_valid_id_o & signal195;
  assign if_id_pipe_reg_we = fetch_valid & id_in_ready_i;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) instr_valid_id_o_t0 <= 1'h0;
    else instr_valid_id_o_t0 <= instr_valid_id_d_t0;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) instr_new_id_o_t0 <= 1'h0;
    else instr_new_id_o_t0 <= if_id_pipe_reg_we_t0;
  assign signal025 = signal192 & pc_set_i;
  assign signal028 = fetch_valid_t0 & signal193;
  assign signal031 = if_id_pipe_reg_we_t0 & signal194;
  assign signal034 = instr_valid_id_o_t0 & signal195;
  assign signal037 = fetch_valid_t0 & id_in_ready_i;
  assign signal026 = pc_set_i_t0 & signal191;
  assign signal029 = fetch_err_t0 & fetch_valid;
  assign signal032 = pc_set_i_t0 & if_id_pipe_reg_we;
  assign signal035 = instr_valid_clear_i_t0 & instr_valid_id_o;
  assign signal038 = id_in_ready_i_t0 & fetch_valid;
  assign signal027 = signal192 & pc_set_i_t0;
  assign signal030 = fetch_valid_t0 & fetch_err_t0;
  assign signal033 = if_id_pipe_reg_we_t0 & pc_set_i_t0;
  assign signal036 = instr_valid_id_o_t0 & instr_valid_clear_i_t0;
  assign signal039 = fetch_valid_t0 & id_in_ready_i_t0;
  assign signal104 = signal025 | signal026;
  assign signal105 = signal028 | signal029;
  assign signal106 = signal031 | signal032;
  assign signal107 = signal034 | signal035;
  assign signal108 = signal037 | signal038;
  assign csr_mtvec_init_o_t0 = signal104 | signal027;
  assign signal001 = signal105 | signal030;
  assign signal003 = signal106 | signal033;
  assign signal005 = signal107 | signal036;
  assign if_id_pipe_reg_we_t0 = signal108 | signal039;
  assign signal161 = pc_if_o ^ pc_id_o;
  assign signal162 = illegal_c_insn ^ illegal_c_insn_id_o;
  assign signal163 = fetch_err_plus2 ^ instr_fetch_err_plus2_o;
  assign signal164 = fetch_rdata[15:0] ^ instr_rdata_c_id_o;
  assign signal165 = fetch_err ^ instr_fetch_err_o;
  assign signal166 = instr_is_compressed ^ instr_is_compressed_id_o;
  assign signal167 = instr_decompressed ^ instr_rdata_alu_id_o;
  assign signal006 = ~ if_id_pipe_reg_we;
  assign signal109 = pc_if_o_t0 | pc_id_o_t0;
  assign signal113 = illegal_c_insn_t0 | illegal_c_insn_id_o_t0;
  assign signal117 = fetch_err_plus2_t0 | instr_fetch_err_plus2_o_t0;
  assign signal121 = fetch_rdata_t0[15:0] | instr_rdata_c_id_o_t0;
  assign signal125 = fetch_err_t0 | instr_fetch_err_o_t0;
  assign signal129 = instr_is_compressed_t0 | instr_is_compressed_id_o_t0;
  assign signal133 = instr_decompressed_t0 | instr_rdata_alu_id_o_t0;
  assign signal110 = signal161 | signal109;
  assign signal114 = signal162 | signal113;
  assign signal118 = signal163 | signal117;
  assign signal122 = signal164 | signal121;
  assign signal126 = signal165 | signal125;
  assign signal130 = signal166 | signal129;
  assign signal134 = signal167 | signal133;
  assign signal040 = { if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we } & pc_if_o_t0;
  assign signal043 = if_id_pipe_reg_we & illegal_c_insn_t0;
  assign signal046 = if_id_pipe_reg_we & fetch_err_plus2_t0;
  assign signal049 = { if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we } & fetch_rdata_t0[15:0];
  assign signal052 = if_id_pipe_reg_we & fetch_err_t0;
  assign signal055 = if_id_pipe_reg_we & instr_is_compressed_t0;
  assign signal058 = { if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we } & instr_decompressed_t0;
  assign signal041 = { signal006, signal006, signal006, signal006, signal006, signal006, signal006, signal006, signal006, signal006, signal006, signal006, signal006, signal006, signal006, signal006, signal006, signal006, signal006, signal006, signal006, signal006, signal006, signal006, signal006, signal006, signal006, signal006, signal006, signal006, signal006, signal006 } & pc_id_o_t0;
  assign signal044 = signal006 & illegal_c_insn_id_o_t0;
  assign signal047 = signal006 & instr_fetch_err_plus2_o_t0;
  assign signal050 = { signal006, signal006, signal006, signal006, signal006, signal006, signal006, signal006, signal006, signal006, signal006, signal006, signal006, signal006, signal006, signal006 } & instr_rdata_c_id_o_t0;
  assign signal053 = signal006 & instr_fetch_err_o_t0;
  assign signal056 = signal006 & instr_is_compressed_id_o_t0;
  assign signal059 = { signal006, signal006, signal006, signal006, signal006, signal006, signal006, signal006, signal006, signal006, signal006, signal006, signal006, signal006, signal006, signal006, signal006, signal006, signal006, signal006, signal006, signal006, signal006, signal006, signal006, signal006, signal006, signal006, signal006, signal006, signal006, signal006 } & instr_rdata_alu_id_o_t0;
  assign signal042 = signal110 & if_id_pipe_reg_we_t0;
  assign signal045 = signal114 & if_id_pipe_reg_we_t0;
  assign signal048 = signal118 & if_id_pipe_reg_we_t0;
  assign signal051 = signal122 & if_id_pipe_reg_we_t0;
  assign signal054 = signal126 & if_id_pipe_reg_we_t0;
  assign signal057 = signal130 & if_id_pipe_reg_we_t0;
  assign signal060 = signal134 & if_id_pipe_reg_we_t0;
  assign signal111 = signal040 | signal041;
  assign signal115 = signal043 | signal044;
  assign signal119 = signal046 | signal047;
  assign signal123 = signal049 | signal050;
  assign signal127 = signal052 | signal053;
  assign signal131 = signal055 | signal056;
  assign signal135 = signal058 | signal059;
  assign signal112 = signal111 | signal042;
  assign signal116 = signal115 | signal045;
  assign signal120 = signal119 | signal048;
  assign signal124 = signal123 | signal051;
  assign signal128 = signal127 | signal054;
  assign signal132 = signal131 | signal057;
  assign signal136 = signal135 | signal060;
  always_ff @(posedge clk_i)
    pc_id_o_t0 <= signal112;
  always_ff @(posedge clk_i)
    illegal_c_insn_id_o_t0 <= signal116;
  always_ff @(posedge clk_i)
    instr_fetch_err_plus2_o_t0 <= signal120;
  always_ff @(posedge clk_i)
    instr_rdata_c_id_o_t0 <= signal124;
  always_ff @(posedge clk_i)
    instr_fetch_err_o_t0 <= signal128;
  always_ff @(posedge clk_i)
    instr_is_compressed_id_o_t0 <= signal132;
  always_ff @(posedge clk_i)
    instr_rdata_alu_id_o_t0 <= signal136;
  assign signal022 = | pc_mux_i_t0;
  assign signal023 = | exc_pc_mux_i_t0;
  assign signal018 = ~ pc_mux_i_t0;
  assign signal021 = ~ exc_pc_mux_i_t0;
  assign signal088 = pc_mux_i & signal018;
  assign signal096 = exc_pc_mux_i & signal021;
  assign signal092 = 3'h4 & signal018;
  assign signal093 = 3'h3 & signal018;
  assign signal094 = 3'h2 & signal018;
  assign signal095 = 3'h1 & signal018;
  assign signal097 = 2'h3 & signal021;
  assign signal098 = 2'h2 & signal021;
  assign signal099 = 2'h1 & signal021;
  assign signal174 = signal088 == signal092;
  assign signal175 = signal088 == signal093;
  assign signal176 = signal088 == signal094;
  assign signal177 = signal088 == signal095;
  assign signal178 = signal096 == signal097;
  assign signal179 = signal096 == signal098;
  assign signal180 = signal096 == signal099;
  assign signal197 = signal174 & signal022;
  assign signal199 = signal175 & signal022;
  assign signal201 = signal176 & signal022;
  assign signal203 = signal177 & signal022;
  assign signal205 = signal178 & signal023;
  assign signal207 = signal179 & signal023;
  assign signal209 = signal180 & signal023;
  always_ff @(posedge clk_i)
    if (if_id_pipe_reg_we) pc_id_o <= pc_if_o;
  always_ff @(posedge clk_i)
    if (if_id_pipe_reg_we) illegal_c_insn_id_o <= illegal_c_insn;
  always_ff @(posedge clk_i)
    if (if_id_pipe_reg_we) instr_fetch_err_plus2_o <= fetch_err_plus2;
  always_ff @(posedge clk_i)
    if (if_id_pipe_reg_we) instr_rdata_c_id_o <= fetch_rdata[15:0];
  always_ff @(posedge clk_i)
    if (if_id_pipe_reg_we) instr_fetch_err_o <= fetch_err;
  always_ff @(posedge clk_i)
    if (if_id_pipe_reg_we) instr_is_compressed_id_o <= instr_is_compressed;
  always_ff @(posedge clk_i)
    if (if_id_pipe_reg_we) instr_rdata_alu_id_o <= instr_decompressed;
  assign signal024 = ! signal088;
  assign signal192 = signal024 & signal022;
  assign signal011 = ~ { signal196, signal196, signal196, signal196, signal196, signal196, signal196, signal196, signal196, signal196, signal196, signal196, signal196, signal196, signal196, signal196, signal196, signal196, signal196, signal196, signal196, signal196, signal196, signal196, signal196, signal196, signal196, signal196, signal196, signal196, signal196, signal196 };
  assign signal012 = ~ { signal202, signal202, signal202, signal202, signal202, signal202, signal202, signal202, signal202, signal202, signal202, signal202, signal202, signal202, signal202, signal202, signal202, signal202, signal202, signal202, signal202, signal202, signal202, signal202, signal202, signal202, signal202, signal202, signal202, signal202, signal202, signal202 };
  assign signal013 = ~ { signal200, signal200, signal200, signal200, signal200, signal200, signal200, signal200, signal200, signal200, signal200, signal200, signal200, signal200, signal200, signal200, signal200, signal200, signal200, signal200, signal200, signal200, signal200, signal200, signal200, signal200, signal200, signal200, signal200, signal200, signal200, signal200 };
  assign signal014 = ~ { signal100, signal100, signal100, signal100, signal100, signal100, signal100, signal100, signal100, signal100, signal100, signal100, signal100, signal100, signal100, signal100, signal100, signal100, signal100, signal100, signal100, signal100, signal100, signal100, signal100, signal100, signal100, signal100, signal100, signal100, signal100, signal100 };
  assign signal015 = ~ { signal204, signal204, signal204, signal204, signal204, signal204, signal204, signal204, signal204, signal204, signal204, signal204, signal204, signal204, signal204, signal204, signal204, signal204, signal204, signal204, signal204, signal204, signal204, signal204, signal204, signal204, signal204, signal204, signal204, signal204, signal204, signal204 };
  assign signal016 = ~ { signal208, signal208, signal208, signal208, signal208, signal208, signal208, signal208, signal208, signal208, signal208, signal208, signal208, signal208, signal208, signal208, signal208, signal208, signal208, signal208, signal208, signal208, signal208, signal208, signal208, signal208, signal208, signal208, signal208, signal208, signal208, signal208 };
  assign signal017 = ~ { signal102, signal102, signal102, signal102, signal102, signal102, signal102, signal102, signal102, signal102, signal102, signal102, signal102, signal102, signal102, signal102, signal102, signal102, signal102, signal102, signal102, signal102, signal102, signal102, signal102, signal102, signal102, signal102, signal102, signal102, signal102, signal102 };
  assign signal139 = { signal197, signal197, signal197, signal197, signal197, signal197, signal197, signal197, signal197, signal197, signal197, signal197, signal197, signal197, signal197, signal197, signal197, signal197, signal197, signal197, signal197, signal197, signal197, signal197, signal197, signal197, signal197, signal197, signal197, signal197, signal197, signal197 } | signal011;
  assign signal142 = { signal203, signal203, signal203, signal203, signal203, signal203, signal203, signal203, signal203, signal203, signal203, signal203, signal203, signal203, signal203, signal203, signal203, signal203, signal203, signal203, signal203, signal203, signal203, signal203, signal203, signal203, signal203, signal203, signal203, signal203, signal203, signal203 } | signal012;
  assign signal145 = { signal201, signal201, signal201, signal201, signal201, signal201, signal201, signal201, signal201, signal201, signal201, signal201, signal201, signal201, signal201, signal201, signal201, signal201, signal201, signal201, signal201, signal201, signal201, signal201, signal201, signal201, signal201, signal201, signal201, signal201, signal201, signal201 } | signal013;
  assign signal148 = { signal101, signal101, signal101, signal101, signal101, signal101, signal101, signal101, signal101, signal101, signal101, signal101, signal101, signal101, signal101, signal101, signal101, signal101, signal101, signal101, signal101, signal101, signal101, signal101, signal101, signal101, signal101, signal101, signal101, signal101, signal101, signal101 } | signal014;
  assign signal151 = { signal205, signal205, signal205, signal205, signal205, signal205, signal205, signal205, signal205, signal205, signal205, signal205, signal205, signal205, signal205, signal205, signal205, signal205, signal205, signal205, signal205, signal205, signal205, signal205, signal205, signal205, signal205, signal205, signal205, signal205, signal205, signal205 } | signal015;
  assign signal154 = { signal209, signal209, signal209, signal209, signal209, signal209, signal209, signal209, signal209, signal209, signal209, signal209, signal209, signal209, signal209, signal209, signal209, signal209, signal209, signal209, signal209, signal209, signal209, signal209, signal209, signal209, signal209, signal209, signal209, signal209, signal209, signal209 } | signal016;
  assign signal157 = { signal103, signal103, signal103, signal103, signal103, signal103, signal103, signal103, signal103, signal103, signal103, signal103, signal103, signal103, signal103, signal103, signal103, signal103, signal103, signal103, signal103, signal103, signal103, signal103, signal103, signal103, signal103, signal103, signal103, signal103, signal103, signal103 } | signal017;
  assign signal140 = { signal197, signal197, signal197, signal197, signal197, signal197, signal197, signal197, signal197, signal197, signal197, signal197, signal197, signal197, signal197, signal197, signal197, signal197, signal197, signal197, signal197, signal197, signal197, signal197, signal197, signal197, signal197, signal197, signal197, signal197, signal197, signal197 } | { signal196, signal196, signal196, signal196, signal196, signal196, signal196, signal196, signal196, signal196, signal196, signal196, signal196, signal196, signal196, signal196, signal196, signal196, signal196, signal196, signal196, signal196, signal196, signal196, signal196, signal196, signal196, signal196, signal196, signal196, signal196, signal196 };
  assign signal143 = { signal203, signal203, signal203, signal203, signal203, signal203, signal203, signal203, signal203, signal203, signal203, signal203, signal203, signal203, signal203, signal203, signal203, signal203, signal203, signal203, signal203, signal203, signal203, signal203, signal203, signal203, signal203, signal203, signal203, signal203, signal203, signal203 } | { signal202, signal202, signal202, signal202, signal202, signal202, signal202, signal202, signal202, signal202, signal202, signal202, signal202, signal202, signal202, signal202, signal202, signal202, signal202, signal202, signal202, signal202, signal202, signal202, signal202, signal202, signal202, signal202, signal202, signal202, signal202, signal202 };
  assign signal146 = { signal201, signal201, signal201, signal201, signal201, signal201, signal201, signal201, signal201, signal201, signal201, signal201, signal201, signal201, signal201, signal201, signal201, signal201, signal201, signal201, signal201, signal201, signal201, signal201, signal201, signal201, signal201, signal201, signal201, signal201, signal201, signal201 } | { signal200, signal200, signal200, signal200, signal200, signal200, signal200, signal200, signal200, signal200, signal200, signal200, signal200, signal200, signal200, signal200, signal200, signal200, signal200, signal200, signal200, signal200, signal200, signal200, signal200, signal200, signal200, signal200, signal200, signal200, signal200, signal200 };
  assign signal149 = { signal101, signal101, signal101, signal101, signal101, signal101, signal101, signal101, signal101, signal101, signal101, signal101, signal101, signal101, signal101, signal101, signal101, signal101, signal101, signal101, signal101, signal101, signal101, signal101, signal101, signal101, signal101, signal101, signal101, signal101, signal101, signal101 } | { signal100, signal100, signal100, signal100, signal100, signal100, signal100, signal100, signal100, signal100, signal100, signal100, signal100, signal100, signal100, signal100, signal100, signal100, signal100, signal100, signal100, signal100, signal100, signal100, signal100, signal100, signal100, signal100, signal100, signal100, signal100, signal100 };
  assign signal152 = { signal205, signal205, signal205, signal205, signal205, signal205, signal205, signal205, signal205, signal205, signal205, signal205, signal205, signal205, signal205, signal205, signal205, signal205, signal205, signal205, signal205, signal205, signal205, signal205, signal205, signal205, signal205, signal205, signal205, signal205, signal205, signal205 } | { signal204, signal204, signal204, signal204, signal204, signal204, signal204, signal204, signal204, signal204, signal204, signal204, signal204, signal204, signal204, signal204, signal204, signal204, signal204, signal204, signal204, signal204, signal204, signal204, signal204, signal204, signal204, signal204, signal204, signal204, signal204, signal204 };
  assign signal155 = { signal209, signal209, signal209, signal209, signal209, signal209, signal209, signal209, signal209, signal209, signal209, signal209, signal209, signal209, signal209, signal209, signal209, signal209, signal209, signal209, signal209, signal209, signal209, signal209, signal209, signal209, signal209, signal209, signal209, signal209, signal209, signal209 } | { signal208, signal208, signal208, signal208, signal208, signal208, signal208, signal208, signal208, signal208, signal208, signal208, signal208, signal208, signal208, signal208, signal208, signal208, signal208, signal208, signal208, signal208, signal208, signal208, signal208, signal208, signal208, signal208, signal208, signal208, signal208, signal208 };
  assign signal158 = { signal103, signal103, signal103, signal103, signal103, signal103, signal103, signal103, signal103, signal103, signal103, signal103, signal103, signal103, signal103, signal103, signal103, signal103, signal103, signal103, signal103, signal103, signal103, signal103, signal103, signal103, signal103, signal103, signal103, signal103, signal103, signal103 } | { signal102, signal102, signal102, signal102, signal102, signal102, signal102, signal102, signal102, signal102, signal102, signal102, signal102, signal102, signal102, signal102, signal102, signal102, signal102, signal102, signal102, signal102, signal102, signal102, signal102, signal102, signal102, signal102, signal102, signal102, signal102, signal102 };
  assign signal067 = csr_mepc_i_t0 & signal139;
  assign signal070 = { boot_addr_i_t0[31:8], 8'h00 } & signal142;
  assign signal073 = signal184 & signal145;
  assign signal076 = signal186 & signal148;
  assign signal079 = 32'd0 & signal151;
  assign signal082 = { csr_mtvec_i_t0[31:8], 8'h00 } & signal154;
  assign signal085 = signal190 & signal157;
  assign signal068 = csr_depc_i_t0 & signal140;
  assign signal071 = branch_target_ex_i_t0 & signal143;
  assign signal074 = exc_pc_t0 & signal146;
  assign signal077 = signal182 & signal149;
  assign signal080 = 32'd0 & signal152;
  assign signal083 = { csr_mtvec_i_t0[31:8], 1'h0, exc_cause_t0[4:0], 2'h0 } & signal155;
  assign signal086 = signal188 & signal158;
  assign signal141 = signal067 | signal068;
  assign signal144 = signal070 | signal071;
  assign signal147 = signal073 | signal074;
  assign signal150 = signal076 | signal077;
  assign signal153 = signal079 | signal080;
  assign signal156 = signal082 | signal083;
  assign signal159 = signal085 | signal086;
  assign signal168 = csr_mepc_i ^ csr_depc_i;
  assign signal169 = { boot_addr_i[31:8], 8'h80 } ^ branch_target_ex_i;
  assign signal170 = signal183 ^ exc_pc;
  assign signal171 = signal185 ^ signal181;
  assign signal172 = { csr_mtvec_i[31:8], 8'h00 } ^ { csr_mtvec_i[31:8], 1'h0, exc_cause[4:0], 2'h0 };
  assign signal173 = signal189 ^ signal187;
  assign signal069 = { signal197, signal197, signal197, signal197, signal197, signal197, signal197, signal197, signal197, signal197, signal197, signal197, signal197, signal197, signal197, signal197, signal197, signal197, signal197, signal197, signal197, signal197, signal197, signal197, signal197, signal197, signal197, signal197, signal197, signal197, signal197, signal197 } & signal168;
  assign signal072 = { signal203, signal203, signal203, signal203, signal203, signal203, signal203, signal203, signal203, signal203, signal203, signal203, signal203, signal203, signal203, signal203, signal203, signal203, signal203, signal203, signal203, signal203, signal203, signal203, signal203, signal203, signal203, signal203, signal203, signal203, signal203, signal203 } & signal169;
  assign signal075 = { signal201, signal201, signal201, signal201, signal201, signal201, signal201, signal201, signal201, signal201, signal201, signal201, signal201, signal201, signal201, signal201, signal201, signal201, signal201, signal201, signal201, signal201, signal201, signal201, signal201, signal201, signal201, signal201, signal201, signal201, signal201, signal201 } & signal170;
  assign signal078 = { signal101, signal101, signal101, signal101, signal101, signal101, signal101, signal101, signal101, signal101, signal101, signal101, signal101, signal101, signal101, signal101, signal101, signal101, signal101, signal101, signal101, signal101, signal101, signal101, signal101, signal101, signal101, signal101, signal101, signal101, signal101, signal101 } & signal171;
  assign signal081 = { signal205, signal205, signal205, signal205, signal205, signal205, signal205, signal205, signal205, signal205, signal205, signal205, signal205, signal205, signal205, signal205, signal205, signal205, signal205, signal205, signal205, signal205, signal205, signal205, signal205, signal205, signal205, signal205, signal205, signal205, signal205, signal205 } & 32'd8;
  assign signal084 = { signal209, signal209, signal209, signal209, signal209, signal209, signal209, signal209, signal209, signal209, signal209, signal209, signal209, signal209, signal209, signal209, signal209, signal209, signal209, signal209, signal209, signal209, signal209, signal209, signal209, signal209, signal209, signal209, signal209, signal209, signal209, signal209 } & signal172;
  assign signal087 = { signal103, signal103, signal103, signal103, signal103, signal103, signal103, signal103, signal103, signal103, signal103, signal103, signal103, signal103, signal103, signal103, signal103, signal103, signal103, signal103, signal103, signal103, signal103, signal103, signal103, signal103, signal103, signal103, signal103, signal103, signal103, signal103 } & signal173;
  assign signal182 = signal069 | signal141;
  assign signal184 = signal072 | signal144;
  assign signal186 = signal075 | signal147;
  assign fetch_addr_n_t0 = signal078 | signal150;
  assign signal188 = signal081 | signal153;
  assign signal190 = signal084 | signal156;
  assign exc_pc_t0 = signal087 | signal159;
  assign signal007 = ~ signal198;
  assign signal009 = ~ signal206;
  assign signal019 = ~ signal002;
  assign signal008 = ~ signal196;
  assign signal010 = ~ signal204;
  assign signal020 = ~ signal004;
  assign signal061 = signal199 & signal008;
  assign signal064 = signal207 & signal010;
  assign signal089 = signal003 & signal020;
  assign signal062 = signal197 & signal007;
  assign signal065 = signal205 & signal009;
  assign signal090 = signal005 & signal019;
  assign signal063 = signal199 & signal197;
  assign signal066 = signal207 & signal205;
  assign signal091 = signal003 & signal005;
  assign signal137 = signal061 | signal062;
  assign signal138 = signal064 | signal065;
  assign signal160 = signal089 | signal090;
  assign signal101 = signal137 | signal063;
  assign signal103 = signal138 | signal066;
  assign instr_valid_id_d_t0 = signal160 | signal091;
  assign signal100 = signal198 | signal196;
  assign signal102 = signal206 | signal204;
  assign signal181 = signal196 ? csr_depc_i : csr_mepc_i;
  assign signal183 = signal202 ? branch_target_ex_i : { boot_addr_i[31:8], 8'h80 };
  assign signal185 = signal200 ? exc_pc : signal183;
  assign fetch_addr_n = signal100 ? signal181 : signal185;
  assign signal187 = signal204 ? 32'd437323784 : 32'd437323776;
  assign signal189 = signal208 ? { csr_mtvec_i[31:8], 1'h0, exc_cause[4:0], 2'h0 } : { csr_mtvec_i[31:8], 8'h00 };
  assign exc_pc = signal102 ? signal187 : signal189;
  assign signal191 = ! pc_mux_i;
  assign signal193 = ~ fetch_err;
  assign signal194 = ~ pc_set_i;
  assign signal195 = ~ instr_valid_clear_i;
  assign instr_valid_id_d = signal002 | signal004;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) instr_valid_id_o <= 1'h0;
    else instr_valid_id_o <= instr_valid_id_d;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) instr_new_id_o <= 1'h0;
    else instr_new_id_o <= if_id_pipe_reg_we;
  assign signal196 = pc_mux_i == 3'h4;
  assign signal198 = pc_mux_i == 3'h3;
  assign signal200 = pc_mux_i == 3'h2;
  assign signal202 = pc_mux_i == 3'h1;
  assign signal204 = exc_pc_mux_i == 2'h3;
  assign signal206 = exc_pc_mux_i == 2'h2;
  assign signal208 = exc_pc_mux_i == 2'h1;
  auxy_ibex_compressed_decoder compressed_decoder_i (
    .clk_i(clk_i),
    .illegal_instr_o(illegal_c_insn),
    .illegal_instr_o_t0(illegal_c_insn_t0),
    .instr_i(fetch_rdata),
    .instr_i_t0(fetch_rdata_t0),
    .instr_o(instr_decompressed),
    .instr_o_t0(instr_decompressed_t0),
    .is_compressed_o(instr_is_compressed),
    .is_compressed_o_t0(instr_is_compressed_t0),
    .rst_ni(rst_ni),
    .valid_i(signal000),
    .valid_i_t0(signal001)
  );
  paramodauxy_ibex_prefetch_bufferBranchPredictor10  \gen_prefetch_buffer.prefetch_buffer_i  (
    .addr_i({ fetch_addr_n[31:1], 1'h0 }),
    .addr_i_t0({ fetch_addr_n_t0[31:1], 1'h0 }),
    .addr_o(pc_if_o),
    .addr_o_t0(pc_if_o_t0),
    .branch_i(pc_set_i),
    .branch_i_t0(pc_set_i_t0),
    .branch_mispredict_i(nt_branch_mispredict_i),
    .branch_mispredict_i_t0(nt_branch_mispredict_i_t0),
    .branch_spec_i(pc_set_spec_i),
    .branch_spec_i_t0(pc_set_spec_i_t0),
    .busy_o(if_busy_o),
    .busy_o_t0(if_busy_o_t0),
    .clk_i(clk_i),
    .err_o(fetch_err),
    .err_o_t0(fetch_err_t0),
    .err_plus2_o(fetch_err_plus2),
    .err_plus2_o_t0(fetch_err_plus2_t0),
    .instr_addr_o(instr_addr_o),
    .instr_addr_o_t0(instr_addr_o_t0),
    .instr_err_i(instr_err_i),
    .instr_err_i_t0(instr_err_i_t0),
    .instr_gnt_i(instr_gnt_i),
    .instr_gnt_i_t0(instr_gnt_i_t0),
    .instr_pmp_err_i(instr_pmp_err_i),
    .instr_pmp_err_i_t0(instr_pmp_err_i_t0),
    .instr_rdata_i(instr_rdata_i),
    .instr_rdata_i_t0(instr_rdata_i_t0),
    .instr_req_o(instr_req_o),
    .instr_req_o_t0(instr_req_o_t0),
    .instr_rvalid_i(instr_rvalid_i),
    .instr_rvalid_i_t0(instr_rvalid_i_t0),
    .predicted_branch_i(1'h0),
    .predicted_branch_i_t0(1'h0),
    .rdata_o(fetch_rdata),
    .rdata_o_t0(fetch_rdata_t0),
    .ready_i(id_in_ready_i),
    .ready_i_t0(id_in_ready_i_t0),
    .req_i(req_i),
    .req_i_t0(req_i_t0),
    .rst_ni(rst_ni),
    .valid_o(fetch_valid),
    .valid_o_t0(fetch_valid_t0)
  );
  assign dummy_instr_id_o = 1'h0;
  assign dummy_instr_id_o_t0 = 1'h0;
  assign ic_data_addr_o = 8'h00;
  assign ic_data_addr_o_t0 = 8'h00;
  assign ic_data_req_o = 2'h0;
  assign ic_data_req_o_t0 = 2'h0;
  assign ic_data_wdata_o = 64'h0000000000000000;
  assign ic_data_wdata_o_t0 = 64'h0000000000000000;
  assign ic_data_write_o = 1'h0;
  assign ic_data_write_o_t0 = 1'h0;
  assign ic_tag_addr_o = 8'h00;
  assign ic_tag_addr_o_t0 = 8'h00;
  assign ic_tag_req_o = 2'h0;
  assign ic_tag_req_o_t0 = 2'h0;
  assign ic_tag_wdata_o = 22'h000000;
  assign ic_tag_wdata_o_t0 = 22'h000000;
  assign ic_tag_write_o = 1'h0;
  assign ic_tag_write_o_t0 = 1'h0;
  assign instr_bp_taken_o = 1'h0;
  assign instr_bp_taken_o_t0 = 1'h0;
  assign instr_rdata_id_o = instr_rdata_alu_id_o;
  assign instr_rdata_id_o_t0 = instr_rdata_alu_id_o_t0;
  assign pc_mismatch_alert_o = 1'h0;
  assign pc_mismatch_alert_o_t0 = 1'h0;
endmodule

module paramod2736aa8a03348385795fda019fbdaaafd7f2ecf9auxy_ibex_csr (clk_i, rst_ni, wr_data_i, wr_en_i, rd_data_o, rd_error_o, rd_data_o_t0, rd_error_o_t0, wr_data_i_t0, wr_en_i_t0);
  wire _00_;
  wire [5:0] _01_;
  wire [5:0] _02_;
  wire [5:0] _03_;
  wire [5:0] _04_;
  wire [5:0] _05_;
  wire [5:0] _06_;
  wire [5:0] _07_;
  wire [5:0] _08_;
  input clk_i;
  wire clk_i;
  output [5:0] rd_data_o;
  reg [5:0] rd_data_o;
  output [5:0] rd_data_o_t0;
  reg [5:0] rd_data_o_t0;
  output rd_error_o;
  wire rd_error_o;
  output rd_error_o_t0;
  wire rd_error_o_t0;
  input rst_ni;
  wire rst_ni;
  input [5:0] wr_data_i;
  wire [5:0] wr_data_i;
  input [5:0] wr_data_i_t0;
  wire [5:0] wr_data_i_t0;
  input wr_en_i;
  wire wr_en_i;
  input wr_en_i_t0;
  wire wr_en_i_t0;
  assign _00_ = ~ wr_en_i;
  assign _08_ = wr_data_i ^ rd_data_o;
  assign _04_ = wr_data_i_t0 | rd_data_o_t0;
  assign _05_ = _08_ | _04_;
  assign _01_ = { wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i } & wr_data_i_t0;
  assign _02_ = { _00_, _00_, _00_, _00_, _00_, _00_ } & rd_data_o_t0;
  assign _03_ = _05_ & { wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0 };
  assign _06_ = _01_ | _02_;
  assign _07_ = _06_ | _03_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) rd_data_o_t0 <= 6'h00;
    else rd_data_o_t0 <= _07_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) rd_data_o <= 6'h00;
    else if (wr_en_i) rd_data_o <= wr_data_i;
  assign rd_error_o = 1'h0;
  assign rd_error_o_t0 = 1'h0;
endmodule

module paramod4033ffde0d007f439ab68268c14c7a2b914b41b4auxy_prim_fifo_sync (clk_i, rst_ni, clr_i, wvalid_i, wready_o, wdata_i, rvalid_o, rready_i, rdata_o, full_o, depth_o, rready_i_t0, rvalid_o_t0, wdata_i_t0, wready_o_t0, wvalid_i_t0, clr_i_t0, depth_o_t0, full_o_t0, rdata_o_t0);
  input clk_i;
  wire clk_i;
  input clr_i;
  wire clr_i;
  input clr_i_t0;
  wire clr_i_t0;
  output depth_o;
  wire depth_o;
  output depth_o_t0;
  wire depth_o_t0;
  output full_o;
  wire full_o;
  output full_o_t0;
  wire full_o_t0;
  output [64:0] rdata_o;
  wire [64:0] rdata_o;
  output [64:0] rdata_o_t0;
  wire [64:0] rdata_o_t0;
  input rready_i;
  wire rready_i;
  input rready_i_t0;
  wire rready_i_t0;
  input rst_ni;
  wire rst_ni;
  output rvalid_o;
  wire rvalid_o;
  output rvalid_o_t0;
  wire rvalid_o_t0;
  input [64:0] wdata_i;
  wire [64:0] wdata_i;
  input [64:0] wdata_i_t0;
  wire [64:0] wdata_i_t0;
  output wready_o;
  wire wready_o;
  output wready_o_t0;
  wire wready_o_t0;
  input wvalid_i;
  wire wvalid_i;
  input wvalid_i_t0;
  wire wvalid_i_t0;
  assign depth_o = 1'h0;
  assign depth_o_t0 = 1'h0;
  assign full_o = rready_i;
  assign full_o_t0 = rready_i_t0;
  assign rdata_o = wdata_i;
  assign rdata_o_t0 = wdata_i_t0;
  assign rvalid_o = wvalid_i;
  assign rvalid_o_t0 = wvalid_i_t0;
  assign wready_o = rready_i;
  assign wready_o_t0 = rready_i_t0;
endmodule

module paramod410b37fbfbfa994790f1902c150d2be939cadb3bauxy_ibex_csr (clk_i, rst_ni, wr_data_i, wr_en_i, rd_data_o, rd_error_o, rd_data_o_t0, rd_error_o_t0, wr_data_i_t0, wr_en_i_t0);
  wire _00_;
  wire [2:0] _01_;
  wire [2:0] _02_;
  wire [2:0] _03_;
  wire [2:0] _04_;
  wire [2:0] _05_;
  wire [2:0] _06_;
  wire [2:0] _07_;
  wire [2:0] _08_;
  input clk_i;
  wire clk_i;
  output [2:0] rd_data_o;
  reg [2:0] rd_data_o;
  output [2:0] rd_data_o_t0;
  reg [2:0] rd_data_o_t0;
  output rd_error_o;
  wire rd_error_o;
  output rd_error_o_t0;
  wire rd_error_o_t0;
  input rst_ni;
  wire rst_ni;
  input [2:0] wr_data_i;
  wire [2:0] wr_data_i;
  input [2:0] wr_data_i_t0;
  wire [2:0] wr_data_i_t0;
  input wr_en_i;
  wire wr_en_i;
  input wr_en_i_t0;
  wire wr_en_i_t0;
  assign _00_ = ~ wr_en_i;
  assign _08_ = wr_data_i ^ rd_data_o;
  assign _04_ = wr_data_i_t0 | rd_data_o_t0;
  assign _05_ = _08_ | _04_;
  assign _01_ = { wr_en_i, wr_en_i, wr_en_i } & wr_data_i_t0;
  assign _02_ = { _00_, _00_, _00_ } & rd_data_o_t0;
  assign _03_ = _05_ & { wr_en_i_t0, wr_en_i_t0, wr_en_i_t0 };
  assign _06_ = _01_ | _02_;
  assign _07_ = _06_ | _03_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) rd_data_o_t0 <= 3'h0;
    else rd_data_o_t0 <= _07_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) rd_data_o <= 3'h4;
    else if (wr_en_i) rd_data_o <= wr_data_i;
  assign rd_error_o = 1'h0;
  assign rd_error_o_t0 = 1'h0;
endmodule

module paramod4f46e25470a27719ee9ca03cee1a0827eff766f7auxy_ibex_csr (clk_i, rst_ni, wr_data_i, wr_en_i, rd_data_o, rd_error_o, rd_data_o_t0, rd_error_o_t0, wr_data_i_t0, wr_en_i_t0);
  wire _00_;
  wire [31:0] _01_;
  wire [31:0] _02_;
  wire [31:0] _03_;
  wire [31:0] _04_;
  wire [31:0] _05_;
  wire [31:0] _06_;
  wire [31:0] _07_;
  wire [31:0] _08_;
  input clk_i;
  wire clk_i;
  output [31:0] rd_data_o;
  reg [31:0] rd_data_o;
  output [31:0] rd_data_o_t0;
  reg [31:0] rd_data_o_t0;
  output rd_error_o;
  wire rd_error_o;
  output rd_error_o_t0;
  wire rd_error_o_t0;
  input rst_ni;
  wire rst_ni;
  input [31:0] wr_data_i;
  wire [31:0] wr_data_i;
  input [31:0] wr_data_i_t0;
  wire [31:0] wr_data_i_t0;
  input wr_en_i;
  wire wr_en_i;
  input wr_en_i_t0;
  wire wr_en_i_t0;
  assign _00_ = ~ wr_en_i;
  assign _08_ = wr_data_i ^ rd_data_o;
  assign _04_ = wr_data_i_t0 | rd_data_o_t0;
  assign _05_ = _08_ | _04_;
  assign _01_ = { wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i } & wr_data_i_t0;
  assign _02_ = { _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_ } & rd_data_o_t0;
  assign _03_ = _05_ & { wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0 };
  assign _06_ = _01_ | _02_;
  assign _07_ = _06_ | _03_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) rd_data_o_t0 <= 32'd0;
    else rd_data_o_t0 <= _07_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) rd_data_o <= 32'd1;
    else if (wr_en_i) rd_data_o <= wr_data_i;
  assign rd_error_o = 1'h0;
  assign rd_error_o_t0 = 1'h0;
endmodule

module paramod5714e31d82f2b8816750797f158ebea69a089104auxy_ibex_csr (clk_i, rst_ni, wr_data_i, wr_en_i, rd_data_o, rd_error_o, rd_data_o_t0, rd_error_o_t0, wr_data_i_t0, wr_en_i_t0);
  wire _00_;
  wire [5:0] _01_;
  wire [5:0] _02_;
  wire [5:0] _03_;
  wire [5:0] _04_;
  wire [5:0] _05_;
  wire [5:0] _06_;
  wire [5:0] _07_;
  wire [5:0] _08_;
  input clk_i;
  wire clk_i;
  output [5:0] rd_data_o;
  reg [5:0] rd_data_o;
  output [5:0] rd_data_o_t0;
  reg [5:0] rd_data_o_t0;
  output rd_error_o;
  wire rd_error_o;
  output rd_error_o_t0;
  wire rd_error_o_t0;
  input rst_ni;
  wire rst_ni;
  input [5:0] wr_data_i;
  wire [5:0] wr_data_i;
  input [5:0] wr_data_i_t0;
  wire [5:0] wr_data_i_t0;
  input wr_en_i;
  wire wr_en_i;
  input wr_en_i_t0;
  wire wr_en_i_t0;
  assign _00_ = ~ wr_en_i;
  assign _08_ = wr_data_i ^ rd_data_o;
  assign _04_ = wr_data_i_t0 | rd_data_o_t0;
  assign _05_ = _08_ | _04_;
  assign _01_ = { wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i } & wr_data_i_t0;
  assign _02_ = { _00_, _00_, _00_, _00_, _00_, _00_ } & rd_data_o_t0;
  assign _03_ = _05_ & { wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0 };
  assign _06_ = _01_ | _02_;
  assign _07_ = _06_ | _03_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) rd_data_o_t0 <= 6'h00;
    else rd_data_o_t0 <= _07_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) rd_data_o <= 6'h10;
    else if (wr_en_i) rd_data_o <= wr_data_i;
  assign rd_error_o = 1'h0;
  assign rd_error_o_t0 = 1'h0;
endmodule

module paramod6ae18350b51be32fd7406c5aaac3c7582e0e6af0auxy_prim_flop (clk_i, rst_ni, d_i, q_o, q_o_t0, d_i_t0);
  input clk_i;
  wire clk_i;
  input [3:0] d_i;
  wire [3:0] d_i;
  input [3:0] d_i_t0;
  wire [3:0] d_i_t0;
  output [3:0] q_o;
  wire [3:0] q_o;
  output [3:0] q_o_t0;
  wire [3:0] q_o_t0;
  input rst_ni;
  wire rst_ni;
  paramod6ae18350b51be32fd7406c5aaac3c7582e0e6af0auxy_prim_generic_flop  \gen_generic.u_impl_generic  (
    .clk_i(clk_i),
    .d_i(d_i),
    .d_i_t0(d_i_t0),
    .q_o(q_o),
    .q_o_t0(q_o_t0),
    .rst_ni(rst_ni)
  );
endmodule

module paramod6ae18350b51be32fd7406c5aaac3c7582e0e6af0auxy_prim_flop_2sync (clk_i, rst_ni, d_i, q_o, q_o_t0, d_i_t0);
  input clk_i;
  wire clk_i;
  input [3:0] d_i;
  wire [3:0] d_i;
  input [3:0] d_i_t0;
  wire [3:0] d_i_t0;
  output [3:0] q_o;
  wire [3:0] q_o;
  output [3:0] q_o_t0;
  wire [3:0] q_o_t0;
  input rst_ni;
  wire rst_ni;
  paramod6ae18350b51be32fd7406c5aaac3c7582e0e6af0auxy_prim_generic_flop_2sync  \gen_generic.u_impl_generic  (
    .clk_i(clk_i),
    .d_i(d_i),
    .d_i_t0(d_i_t0),
    .q_o(q_o),
    .q_o_t0(q_o_t0),
    .rst_ni(rst_ni)
  );
endmodule

module paramod6ae18350b51be32fd7406c5aaac3c7582e0e6af0auxy_prim_generic_flop (clk_i, rst_ni, d_i, q_o, q_o_t0, d_i_t0);
  input clk_i;
  wire clk_i;
  input [3:0] d_i;
  wire [3:0] d_i;
  input [3:0] d_i_t0;
  wire [3:0] d_i_t0;
  output [3:0] q_o;
  reg [3:0] q_o;
  output [3:0] q_o_t0;
  reg [3:0] q_o_t0;
  input rst_ni;
  wire rst_ni;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) q_o_t0 <= 4'h0;
    else q_o_t0 <= d_i_t0;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) q_o <= 4'h5;
    else q_o <= d_i;
endmodule

module paramod6ae18350b51be32fd7406c5aaac3c7582e0e6af0auxy_prim_generic_flop_2sync (clk_i, rst_ni, d_i, q_o, q_o_t0, d_i_t0);
  input clk_i;
  wire clk_i;
  input [3:0] d_i;
  wire [3:0] d_i;
  input [3:0] d_i_t0;
  wire [3:0] d_i_t0;
  wire [3:0] intq;
  wire [3:0] intq_t0;
  output [3:0] q_o;
  wire [3:0] q_o;
  output [3:0] q_o_t0;
  wire [3:0] q_o_t0;
  input rst_ni;
  wire rst_ni;
  paramod6ae18350b51be32fd7406c5aaac3c7582e0e6af0auxy_prim_flop  u_sync_1 (
    .clk_i(clk_i),
    .d_i(d_i),
    .d_i_t0(d_i_t0),
    .q_o(intq),
    .q_o_t0(intq_t0),
    .rst_ni(rst_ni)
  );
  paramod6ae18350b51be32fd7406c5aaac3c7582e0e6af0auxy_prim_flop  u_sync_2 (
    .clk_i(clk_i),
    .d_i(intq),
    .d_i_t0(intq_t0),
    .q_o(q_o),
    .q_o_t0(q_o_t0),
    .rst_ni(rst_ni)
  );
endmodule

module paramod85ba01ab5a28334786aba5877c1fe04472f39fbaauxy_ibex_csr (clk_i, rst_ni, wr_data_i, wr_en_i, rd_data_o, rd_error_o, rd_data_o_t0, rd_error_o_t0, wr_data_i_t0, wr_en_i_t0);
  wire _00_;
  wire [31:0] _01_;
  wire [31:0] _02_;
  wire [31:0] _03_;
  wire [31:0] _04_;
  wire [31:0] _05_;
  wire [31:0] _06_;
  wire [31:0] _07_;
  wire [31:0] _08_;
  input clk_i;
  wire clk_i;
  output [31:0] rd_data_o;
  reg [31:0] rd_data_o;
  output [31:0] rd_data_o_t0;
  reg [31:0] rd_data_o_t0;
  output rd_error_o;
  wire rd_error_o;
  output rd_error_o_t0;
  wire rd_error_o_t0;
  input rst_ni;
  wire rst_ni;
  input [31:0] wr_data_i;
  wire [31:0] wr_data_i;
  input [31:0] wr_data_i_t0;
  wire [31:0] wr_data_i_t0;
  input wr_en_i;
  wire wr_en_i;
  input wr_en_i_t0;
  wire wr_en_i_t0;
  assign _00_ = ~ wr_en_i;
  assign _08_ = wr_data_i ^ rd_data_o;
  assign _04_ = wr_data_i_t0 | rd_data_o_t0;
  assign _05_ = _08_ | _04_;
  assign _01_ = { wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i } & wr_data_i_t0;
  assign _02_ = { _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_ } & rd_data_o_t0;
  assign _03_ = _05_ & { wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0 };
  assign _06_ = _01_ | _02_;
  assign _07_ = _06_ | _03_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) rd_data_o_t0 <= 32'd0;
    else rd_data_o_t0 <= _07_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) rd_data_o <= 32'd0;
    else if (wr_en_i) rd_data_o <= wr_data_i;
  assign rd_error_o = 1'h0;
  assign rd_error_o_t0 = 1'h0;
endmodule

module paramod877a50dace05ef79dab022285c3f67914151b286auxy_prim_fifo_sync (clk_i, rst_ni, clr_i, wvalid_i, wready_o, wdata_i, rvalid_o, rready_i, rdata_o, full_o, depth_o, rready_i_t0, rvalid_o_t0, wdata_i_t0, wready_o_t0, wvalid_i_t0, clr_i_t0, depth_o_t0, full_o_t0, rdata_o_t0);
  wire [1:0] _000_;
  wire [1:0] _001_;
  wire [1:0] _002_;
  wire [1:0] _003_;
  wire _004_;
  wire _005_;
  wire _006_;
  wire _007_;
  wire [1:0] _008_;
  wire [1:0] _009_;
  wire [1:0] _010_;
  wire [1:0] _011_;
  wire _012_;
  wire _013_;
  wire _014_;
  wire _015_;
  wire _016_;
  wire _017_;
  wire _018_;
  wire _019_;
  wire _020_;
  wire _021_;
  wire [1:0] _022_;
  wire [1:0] _023_;
  wire _024_;
  wire _025_;
  wire _026_;
  wire [1:0] _027_;
  wire [1:0] _028_;
  wire _029_;
  wire [1:0] _030_;
  wire [1:0] _031_;
  wire [1:0] _032_;
  wire [1:0] _033_;
  wire [1:0] _034_;
  wire [1:0] _035_;
  wire _036_;
  wire _037_;
  wire _038_;
  wire _039_;
  wire [31:0] _040_;
  wire _041_;
  wire _042_;
  wire _043_;
  wire _044_;
  wire _045_;
  wire _046_;
  wire _047_;
  wire _048_;
  wire _049_;
  wire [1:0] _050_;
  wire [1:0] _051_;
  wire _052_;
  wire _053_;
  wire _054_;
  wire _055_;
  wire _056_;
  wire _057_;
  wire _058_;
  wire _059_;
  wire _060_;
  wire _061_;
  wire _062_;
  wire _063_;
  wire _064_;
  wire _065_;
  wire _066_;
  wire _067_;
  wire _068_;
  wire _069_;
  wire [1:0] _070_;
  wire [1:0] _071_;
  wire [1:0] _072_;
  wire [4:0] _073_;
  wire [4:0] _074_;
  wire [4:0] _075_;
  wire [1:0] _076_;
  wire [1:0] _077_;
  wire [1:0] _078_;
  wire [1:0] _079_;
  wire [1:0] _080_;
  wire _081_;
  wire _082_;
  wire [1:0] _083_;
  wire [1:0] _084_;
  wire [1:0] _085_;
  wire [1:0] _086_;
  wire [1:0] _087_;
  wire [1:0] _088_;
  wire [1:0] _089_;
  wire [1:0] _090_;
  wire [1:0] _091_;
  wire [1:0] _092_;
  wire [1:0] _093_;
  wire [1:0] _094_;
  wire [1:0] _095_;
  wire [1:0] _096_;
  wire [1:0] _097_;
  wire [1:0] _098_;
  wire [1:0] _099_;
  wire [1:0] _100_;
  wire [1:0] _101_;
  wire [1:0] _102_;
  wire _103_;
  wire _104_;
  wire _105_;
  wire _106_;
  wire _107_;
  wire _108_;
  wire _109_;
  wire _110_;
  wire [31:0] _111_;
  wire [31:0] _112_;
  wire [31:0] _113_;
  wire _114_;
  wire _115_;
  wire _116_;
  wire [1:0] _117_;
  wire [1:0] _118_;
  wire _119_;
  wire _120_;
  wire _121_;
  wire _122_;
  wire _123_;
  wire _124_;
  wire [1:0] _125_;
  wire [1:0] _126_;
  wire [1:0] _127_;
  wire [1:0] _128_;
  wire [4:0] _129_;
  wire [4:0] _130_;
  wire [4:0] _131_;
  wire [4:0] _132_;
  wire [1:0] _133_;
  wire [1:0] _134_;
  wire [1:0] _135_;
  wire [1:0] _136_;
  wire _137_;
  wire [1:0] _138_;
  wire [1:0] _139_;
  wire [1:0] _140_;
  wire [1:0] _141_;
  wire [1:0] _142_;
  wire [1:0] _143_;
  wire [1:0] _144_;
  wire [1:0] _145_;
  wire [1:0] _146_;
  wire [1:0] _147_;
  wire [1:0] _148_;
  wire [1:0] _149_;
  wire [1:0] _150_;
  wire [1:0] _151_;
  wire [1:0] _152_;
  wire [1:0] _153_;
  wire [1:0] _154_;
  wire _155_;
  wire _156_;
  wire _157_;
  wire _158_;
  wire _159_;
  wire _160_;
  wire _161_;
  wire _162_;
  wire [31:0] _163_;
  wire [31:0] _164_;
  wire [31:0] _165_;
  wire _166_;
  wire [1:0] _167_;
  wire [1:0] _168_;
  wire [1:0] _169_;
  wire [4:0] _170_;
  wire [1:0] _171_;
  wire [1:0] _172_;
  wire [1:0] _173_;
  wire [1:0] _174_;
  wire [1:0] _175_;
  wire [1:0] _176_;
  wire [1:0] _177_;
  wire _178_;
  wire _179_;
  wire _180_;
  wire _181_;
  wire _182_;
  wire _183_;
  wire _184_;
  wire [1:0] _185_;
  wire [1:0] _186_;
  wire [1:0] _187_;
  wire [1:0] _188_;
  wire _189_;
  wire _190_;
  wire _191_;
  wire _192_;
  wire _193_;
  wire _194_;
  wire _195_;
  wire _196_;
  wire _197_;
  wire [1:0] _198_;
  wire [1:0] _199_;
  wire [1:0] _200_;
  wire [1:0] _201_;
  wire _202_;
  wire _203_;
  wire _204_;
  wire _205_;
  wire _206_;
  wire _207_;
  wire [31:0] _208_;
  wire [31:0] _209_;
  wire [1:0] _210_;
  input clk_i;
  wire clk_i;
  input clr_i;
  wire clr_i;
  input clr_i_t0;
  wire clr_i_t0;
  output depth_o;
  wire depth_o;
  output depth_o_t0;
  wire depth_o_t0;
  output full_o;
  wire full_o;
  output full_o_t0;
  wire full_o_t0;
  wire \gen_normal_fifo.empty ;
  wire \gen_normal_fifo.empty_t0 ;
  wire \gen_normal_fifo.fifo_incr_rptr ;
  wire \gen_normal_fifo.fifo_incr_rptr_t0 ;
  wire \gen_normal_fifo.fifo_incr_wptr ;
  wire \gen_normal_fifo.fifo_incr_wptr_t0 ;
  reg [1:0] \gen_normal_fifo.fifo_rptr ;
  reg [1:0] \gen_normal_fifo.fifo_rptr_t0 ;
  reg [1:0] \gen_normal_fifo.fifo_wptr ;
  reg [1:0] \gen_normal_fifo.fifo_wptr_t0 ;
  reg [4:0] \gen_normal_fifo.rdata_int ;
  reg [4:0] \gen_normal_fifo.rdata_int_t0 ;
  reg \gen_normal_fifo.under_rst ;
  reg \gen_normal_fifo.under_rst_t0 ;
  output [4:0] rdata_o;
  wire [4:0] rdata_o;
  output [4:0] rdata_o_t0;
  wire [4:0] rdata_o_t0;
  input rready_i;
  wire rready_i;
  input rready_i_t0;
  wire rready_i_t0;
  input rst_ni;
  wire rst_ni;
  output rvalid_o;
  wire rvalid_o;
  output rvalid_o_t0;
  wire rvalid_o_t0;
  input [4:0] wdata_i;
  wire [4:0] wdata_i;
  input [4:0] wdata_i_t0;
  wire [4:0] wdata_i_t0;
  output wready_o;
  wire wready_o;
  output wready_o_t0;
  wire wready_o_t0;
  input wvalid_i;
  wire wvalid_i;
  input wvalid_i_t0;
  wire wvalid_i_t0;
  assign _006_ = _204_ + \gen_normal_fifo.fifo_wptr [0];
  assign _008_ = \gen_normal_fifo.fifo_wptr  + 2'h1;
  assign _010_ = \gen_normal_fifo.fifo_rptr  + 2'h1;
  assign _012_ = wvalid_i & wready_o;
  assign \gen_normal_fifo.fifo_incr_wptr  = _012_ & _036_;
  assign _014_ = rvalid_o & rready_i;
  assign \gen_normal_fifo.fifo_incr_rptr  = _014_ & _036_;
  assign wready_o = _039_ & _036_;
  assign rvalid_o = _195_ & _036_;
  assign _020_ = ~ _205_;
  assign _022_ = ~ \gen_normal_fifo.fifo_wptr_t0 ;
  assign _023_ = ~ \gen_normal_fifo.fifo_rptr_t0 ;
  assign _048_ = _204_ & _020_;
  assign _050_ = \gen_normal_fifo.fifo_wptr  & _022_;
  assign _051_ = \gen_normal_fifo.fifo_rptr  & _023_;
  assign _183_ = _048_ + _049_;
  assign _185_ = _050_ + 2'h1;
  assign _187_ = _051_ + 2'h1;
  assign _114_ = _204_ | _205_;
  assign _117_ = \gen_normal_fifo.fifo_wptr  | \gen_normal_fifo.fifo_wptr_t0 ;
  assign _118_ = \gen_normal_fifo.fifo_rptr  | \gen_normal_fifo.fifo_rptr_t0 ;
  assign _184_ = _114_ + _115_;
  assign _186_ = _117_ + 2'h1;
  assign _188_ = _118_ + 2'h1;
  assign _166_ = _183_ ^ _184_;
  assign _167_ = _185_ ^ _186_;
  assign _168_ = _187_ ^ _188_;
  assign _116_ = _166_ | _205_;
  assign _009_ = _167_ | \gen_normal_fifo.fifo_wptr_t0 ;
  assign _011_ = _168_ | \gen_normal_fifo.fifo_rptr_t0 ;
  assign _007_ = _116_ | \gen_normal_fifo.fifo_wptr_t0 [0];
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) \gen_normal_fifo.under_rst_t0  <= 1'h0;
    else \gen_normal_fifo.under_rst_t0  <= _005_;
  assign _024_ = ~ _016_;
  assign _026_ = ~ _018_;
  assign _169_ = _002_ ^ \gen_normal_fifo.fifo_wptr ;
  assign _171_ = _000_ ^ \gen_normal_fifo.fifo_rptr ;
  assign _125_ = _003_ | \gen_normal_fifo.fifo_wptr_t0 ;
  assign _133_ = _001_ | \gen_normal_fifo.fifo_rptr_t0 ;
  assign _126_ = _169_ | _125_;
  assign _134_ = _171_ | _133_;
  assign _070_ = { _016_, _016_ } & _003_;
  assign _076_ = { _018_, _018_ } & _001_;
  assign _071_ = { _024_, _024_ } & \gen_normal_fifo.fifo_wptr_t0 ;
  assign _077_ = { _026_, _026_ } & \gen_normal_fifo.fifo_rptr_t0 ;
  assign _072_ = _126_ & { _017_, _017_ };
  assign _078_ = _134_ & { _019_, _019_ };
  assign _127_ = _070_ | _071_;
  assign _135_ = _076_ | _077_;
  assign _128_ = _127_ | _072_;
  assign _136_ = _135_ | _078_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) \gen_normal_fifo.fifo_wptr_t0  <= 2'h0;
    else \gen_normal_fifo.fifo_wptr_t0  <= _128_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) \gen_normal_fifo.fifo_rptr_t0  <= 2'h0;
    else \gen_normal_fifo.fifo_rptr_t0  <= _136_;
  assign _052_ = wvalid_i_t0 & wready_o;
  assign _055_ = _013_ & _036_;
  assign _058_ = rvalid_o_t0 & rready_i;
  assign _061_ = _015_ & _036_;
  assign _064_ = full_o_t0 & _036_;
  assign _067_ = \gen_normal_fifo.empty_t0  & _036_;
  assign _053_ = wready_o_t0 & wvalid_i;
  assign _056_ = \gen_normal_fifo.under_rst_t0  & _012_;
  assign _059_ = rready_i_t0 & rvalid_o;
  assign _062_ = \gen_normal_fifo.under_rst_t0  & _014_;
  assign _065_ = \gen_normal_fifo.under_rst_t0  & _039_;
  assign _068_ = \gen_normal_fifo.under_rst_t0  & _195_;
  assign _054_ = wvalid_i_t0 & wready_o_t0;
  assign _057_ = _013_ & \gen_normal_fifo.under_rst_t0 ;
  assign _060_ = rvalid_o_t0 & rready_i_t0;
  assign _063_ = _015_ & \gen_normal_fifo.under_rst_t0 ;
  assign _066_ = full_o_t0 & \gen_normal_fifo.under_rst_t0 ;
  assign _069_ = \gen_normal_fifo.empty_t0  & \gen_normal_fifo.under_rst_t0 ;
  assign _119_ = _052_ | _053_;
  assign _120_ = _055_ | _056_;
  assign _121_ = _058_ | _059_;
  assign _122_ = _061_ | _062_;
  assign _123_ = _064_ | _065_;
  assign _124_ = _067_ | _068_;
  assign _013_ = _119_ | _054_;
  assign \gen_normal_fifo.fifo_incr_wptr_t0  = _120_ | _057_;
  assign _015_ = _121_ | _060_;
  assign \gen_normal_fifo.fifo_incr_rptr_t0  = _122_ | _063_;
  assign wready_o_t0 = _123_ | _066_;
  assign rvalid_o_t0 = _124_ | _069_;
  assign _170_ = wdata_i ^ \gen_normal_fifo.rdata_int ;
  assign _025_ = ~ \gen_normal_fifo.fifo_incr_wptr ;
  assign _129_ = wdata_i_t0 | \gen_normal_fifo.rdata_int_t0 ;
  assign _130_ = _170_ | _129_;
  assign _073_ = { \gen_normal_fifo.fifo_incr_wptr , \gen_normal_fifo.fifo_incr_wptr , \gen_normal_fifo.fifo_incr_wptr , \gen_normal_fifo.fifo_incr_wptr , \gen_normal_fifo.fifo_incr_wptr  } & wdata_i_t0;
  assign _074_ = { _025_, _025_, _025_, _025_, _025_ } & \gen_normal_fifo.rdata_int_t0 ;
  assign _075_ = _130_ & \gen_normal_fifo.fifo_incr_wptr_t0 ;
  assign _131_ = _073_ | _074_;
  assign _132_ = _131_ | _075_;
  always_ff @(posedge clk_i)
    \gen_normal_fifo.rdata_int_t0  <= _132_;
  assign _044_ = | { \gen_normal_fifo.fifo_rptr_t0 [1], \gen_normal_fifo.fifo_wptr_t0 [1] };
  assign _045_ = | { \gen_normal_fifo.fifo_rptr_t0 , \gen_normal_fifo.fifo_wptr_t0  };
  assign _137_ = \gen_normal_fifo.fifo_wptr_t0 [1] | \gen_normal_fifo.fifo_rptr_t0 [1];
  assign _138_ = \gen_normal_fifo.fifo_wptr_t0  | \gen_normal_fifo.fifo_rptr_t0 ;
  assign _029_ = ~ _137_;
  assign _030_ = ~ _138_;
  assign _081_ = \gen_normal_fifo.fifo_wptr [1] & _029_;
  assign _083_ = \gen_normal_fifo.fifo_wptr  & _030_;
  assign _082_ = \gen_normal_fifo.fifo_rptr [1] & _029_;
  assign _084_ = _210_ & _030_;
  assign _085_ = \gen_normal_fifo.fifo_rptr  & _030_;
  assign _180_ = _081_ == _082_;
  assign _181_ = _083_ == _084_;
  assign _182_ = _083_ == _085_;
  assign _194_ = _180_ & _044_;
  assign full_o_t0 = _181_ & _045_;
  assign \gen_normal_fifo.empty_t0  = _182_ & _045_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) \gen_normal_fifo.fifo_wptr  <= 2'h0;
    else if (_016_) \gen_normal_fifo.fifo_wptr  <= _002_;
  always_ff @(posedge clk_i)
    if (\gen_normal_fifo.fifo_incr_wptr ) \gen_normal_fifo.rdata_int  <= wdata_i;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) \gen_normal_fifo.fifo_rptr  <= 2'h0;
    else if (_018_) \gen_normal_fifo.fifo_rptr  <= _000_;
  assign _042_ = | { \gen_normal_fifo.fifo_incr_wptr_t0 , clr_i_t0 };
  assign _043_ = | { \gen_normal_fifo.fifo_incr_rptr_t0 , clr_i_t0 };
  assign _027_ = ~ { \gen_normal_fifo.fifo_incr_wptr_t0 , clr_i_t0 };
  assign _028_ = ~ { \gen_normal_fifo.fifo_incr_rptr_t0 , clr_i_t0 };
  assign _079_ = { \gen_normal_fifo.fifo_incr_wptr , clr_i } & _027_;
  assign _080_ = { \gen_normal_fifo.fifo_incr_rptr , clr_i } & _028_;
  assign _046_ = ! _079_;
  assign _047_ = ! _080_;
  assign _017_ = _046_ & _042_;
  assign _019_ = _047_ & _043_;
  assign _031_ = ~ { \gen_normal_fifo.fifo_rptr [0], \gen_normal_fifo.fifo_rptr [0] };
  assign _032_ = ~ { \gen_normal_fifo.fifo_incr_rptr , \gen_normal_fifo.fifo_incr_rptr  };
  assign _034_ = ~ { \gen_normal_fifo.fifo_wptr [0], \gen_normal_fifo.fifo_wptr [0] };
  assign _035_ = ~ { \gen_normal_fifo.fifo_incr_wptr , \gen_normal_fifo.fifo_incr_wptr  };
  assign _033_ = ~ { clr_i, clr_i };
  assign _036_ = ~ \gen_normal_fifo.under_rst ;
  assign _038_ = ~ _193_;
  assign _039_ = ~ full_o;
  assign _040_ = ~ { \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty  };
  assign _139_ = { \gen_normal_fifo.fifo_rptr_t0 [0], \gen_normal_fifo.fifo_rptr_t0 [0] } | _031_;
  assign _142_ = { \gen_normal_fifo.fifo_incr_rptr_t0 , \gen_normal_fifo.fifo_incr_rptr_t0  } | _032_;
  assign _148_ = { \gen_normal_fifo.fifo_wptr_t0 [0], \gen_normal_fifo.fifo_wptr_t0 [0] } | _034_;
  assign _151_ = { \gen_normal_fifo.fifo_incr_wptr_t0 , \gen_normal_fifo.fifo_incr_wptr_t0  } | _035_;
  assign _145_ = { clr_i_t0, clr_i_t0 } | _033_;
  assign _159_ = _194_ | _038_;
  assign _162_ = full_o_t0 | _039_;
  assign _163_ = { \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0  } | _040_;
  assign _140_ = { \gen_normal_fifo.fifo_rptr_t0 [0], \gen_normal_fifo.fifo_rptr_t0 [0] } | { \gen_normal_fifo.fifo_rptr [0], \gen_normal_fifo.fifo_rptr [0] };
  assign _143_ = { \gen_normal_fifo.fifo_incr_rptr_t0 , \gen_normal_fifo.fifo_incr_rptr_t0  } | { \gen_normal_fifo.fifo_incr_rptr , \gen_normal_fifo.fifo_incr_rptr  };
  assign _149_ = { \gen_normal_fifo.fifo_wptr_t0 [0], \gen_normal_fifo.fifo_wptr_t0 [0] } | { \gen_normal_fifo.fifo_wptr [0], \gen_normal_fifo.fifo_wptr [0] };
  assign _152_ = { \gen_normal_fifo.fifo_incr_wptr_t0 , \gen_normal_fifo.fifo_incr_wptr_t0  } | { \gen_normal_fifo.fifo_incr_wptr , \gen_normal_fifo.fifo_incr_wptr  };
  assign _146_ = { clr_i_t0, clr_i_t0 } | { clr_i, clr_i };
  assign _155_ = \gen_normal_fifo.under_rst_t0  | \gen_normal_fifo.under_rst ;
  assign _160_ = _194_ | _193_;
  assign _164_ = { \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0  } | { \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty  };
  assign _086_ = { \gen_normal_fifo.fifo_rptr_t0 [1], 1'h0 } & _139_;
  assign _089_ = 2'h0 & _142_;
  assign _092_ = _199_ & _145_;
  assign _095_ = { \gen_normal_fifo.fifo_wptr_t0 [1], 1'h0 } & _148_;
  assign _098_ = 2'h0 & _151_;
  assign _101_ = _201_ & _145_;
  assign _106_ = _007_ & _159_;
  assign _109_ = _207_ & _162_;
  assign _111_ = { 27'h0000000, \gen_normal_fifo.rdata_int_t0  } & _163_;
  assign _087_ = _011_ & _140_;
  assign _090_ = _198_ & _143_;
  assign _096_ = _009_ & _149_;
  assign _099_ = _200_ & _152_;
  assign _093_ = 2'h0 & _146_;
  assign _103_ = \gen_normal_fifo.under_rst_t0  & _155_;
  assign _107_ = _203_ & _160_;
  assign _112_ = 32'd0 & _164_;
  assign _141_ = _086_ | _087_;
  assign _144_ = _089_ | _090_;
  assign _147_ = _092_ | _093_;
  assign _150_ = _095_ | _096_;
  assign _153_ = _098_ | _099_;
  assign _154_ = _101_ | _093_;
  assign _161_ = _106_ | _107_;
  assign _165_ = _111_ | _112_;
  assign _172_ = { _197_, 1'h0 } ^ _010_;
  assign _175_ = { _196_, 1'h0 } ^ _008_;
  assign _179_ = _006_ ^ _202_;
  assign _088_ = { \gen_normal_fifo.fifo_rptr_t0 [0], \gen_normal_fifo.fifo_rptr_t0 [0] } & _172_;
  assign _091_ = { \gen_normal_fifo.fifo_incr_rptr_t0 , \gen_normal_fifo.fifo_incr_rptr_t0  } & _173_;
  assign _094_ = { clr_i_t0, clr_i_t0 } & _174_;
  assign _097_ = { \gen_normal_fifo.fifo_wptr_t0 [0], \gen_normal_fifo.fifo_wptr_t0 [0] } & _175_;
  assign _100_ = { \gen_normal_fifo.fifo_incr_wptr_t0 , \gen_normal_fifo.fifo_incr_wptr_t0  } & _176_;
  assign _102_ = { clr_i_t0, clr_i_t0 } & _177_;
  assign _104_ = \gen_normal_fifo.under_rst_t0  & _036_;
  assign _108_ = _194_ & _179_;
  assign _110_ = full_o_t0 & _041_;
  assign _113_ = { \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0  } & { 27'h0000000, \gen_normal_fifo.rdata_int  };
  assign _198_ = _088_ | _141_;
  assign _199_ = _091_ | _144_;
  assign _001_ = _094_ | _147_;
  assign _200_ = _097_ | _150_;
  assign _201_ = _100_ | _153_;
  assign _003_ = _102_ | _154_;
  assign _005_ = _104_ | _103_;
  assign _207_ = _108_ | _161_;
  assign depth_o_t0 = _110_ | _109_;
  assign { _209_[31:5], rdata_o_t0 } = _113_ | _165_;
  assign _016_ = | { \gen_normal_fifo.fifo_incr_wptr , clr_i };
  assign _018_ = | { \gen_normal_fifo.fifo_incr_rptr , clr_i };
  assign _041_ = ~ _206_;
  assign _021_ = ~ \gen_normal_fifo.fifo_wptr_t0 [0];
  assign _037_ = ~ \gen_normal_fifo.fifo_rptr_t0 [0];
  assign _049_ = \gen_normal_fifo.fifo_wptr [0] & _021_;
  assign _105_ = \gen_normal_fifo.fifo_rptr [0] & _037_;
  assign _115_ = \gen_normal_fifo.fifo_wptr [0] | \gen_normal_fifo.fifo_wptr_t0 [0];
  assign _156_ = \gen_normal_fifo.fifo_rptr [0] | \gen_normal_fifo.fifo_rptr_t0 [0];
  assign _189_ = _115_ - _105_;
  assign _191_ = 1'h1 - _105_;
  assign _190_ = _049_ - _156_;
  assign _192_ = 1'h1 - _156_;
  assign _178_ = _189_ ^ _190_;
  assign _158_ = _191_ ^ _192_;
  assign _157_ = _178_ | \gen_normal_fifo.fifo_wptr_t0 [0];
  assign _203_ = _157_ | \gen_normal_fifo.fifo_rptr_t0 [0];
  assign _205_ = _158_ | \gen_normal_fifo.fifo_rptr_t0 [0];
  assign _193_ = \gen_normal_fifo.fifo_wptr [1] == \gen_normal_fifo.fifo_rptr [1];
  assign full_o = \gen_normal_fifo.fifo_wptr  == _210_;
  assign \gen_normal_fifo.empty  = \gen_normal_fifo.fifo_wptr  == \gen_normal_fifo.fifo_rptr ;
  assign _195_ = ~ \gen_normal_fifo.empty ;
  assign _196_ = ~ \gen_normal_fifo.fifo_wptr [1];
  assign _197_ = ~ \gen_normal_fifo.fifo_rptr [1];
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) \gen_normal_fifo.under_rst  <= 1'h1;
    else \gen_normal_fifo.under_rst  <= _004_;
  assign _173_ = \gen_normal_fifo.fifo_rptr [0] ? _010_ : { _197_, 1'h0 };
  assign _174_ = \gen_normal_fifo.fifo_incr_rptr  ? _173_ : 2'hx;
  assign _000_ = clr_i ? 2'h0 : _174_;
  assign _176_ = \gen_normal_fifo.fifo_wptr [0] ? _008_ : { _196_, 1'h0 };
  assign _177_ = \gen_normal_fifo.fifo_incr_wptr  ? _176_ : 2'hx;
  assign _002_ = clr_i ? 2'h0 : _177_;
  assign _004_ = \gen_normal_fifo.under_rst  ? _036_ : 1'h0;
  assign _202_ = \gen_normal_fifo.fifo_wptr [0] - \gen_normal_fifo.fifo_rptr [0];
  assign _204_ = 1'h1 - \gen_normal_fifo.fifo_rptr [0];
  assign _206_ = _193_ ? _202_ : _006_;
  assign depth_o = full_o ? 1'h1 : _206_;
  assign { _208_[31:5], rdata_o } = \gen_normal_fifo.empty  ? 32'd0 : { 27'h0000000, \gen_normal_fifo.rdata_int  };
  assign _210_ = \gen_normal_fifo.fifo_rptr  ^ 2'h2;
  assign _208_[4:0] = rdata_o;
  assign _209_[4:0] = rdata_o_t0;
endmodule

module paramod9a435d8f6db004a67362aa9a56f32ea481a74dbeauxy_ibex_csr (clk_i, rst_ni, wr_data_i, wr_en_i, rd_data_o, rd_error_o, rd_data_o_t0, rd_error_o_t0, wr_data_i_t0, wr_en_i_t0);
  wire _00_;
  wire [31:0] _01_;
  wire [31:0] _02_;
  wire [31:0] _03_;
  wire [31:0] _04_;
  wire [31:0] _05_;
  wire [31:0] _06_;
  wire [31:0] _07_;
  wire [31:0] _08_;
  input clk_i;
  wire clk_i;
  output [31:0] rd_data_o;
  reg [31:0] rd_data_o;
  output [31:0] rd_data_o_t0;
  reg [31:0] rd_data_o_t0;
  output rd_error_o;
  wire rd_error_o;
  output rd_error_o_t0;
  wire rd_error_o_t0;
  input rst_ni;
  wire rst_ni;
  input [31:0] wr_data_i;
  wire [31:0] wr_data_i;
  input [31:0] wr_data_i_t0;
  wire [31:0] wr_data_i_t0;
  input wr_en_i;
  wire wr_en_i;
  input wr_en_i_t0;
  wire wr_en_i_t0;
  assign _00_ = ~ wr_en_i;
  assign _08_ = wr_data_i ^ rd_data_o;
  assign _04_ = wr_data_i_t0 | rd_data_o_t0;
  assign _05_ = _08_ | _04_;
  assign _01_ = { wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i } & wr_data_i_t0;
  assign _02_ = { _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_ } & rd_data_o_t0;
  assign _03_ = _05_ & { wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0 };
  assign _06_ = _01_ | _02_;
  assign _07_ = _06_ | _03_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) rd_data_o_t0 <= 32'd0;
    else rd_data_o_t0 <= _07_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) rd_data_o <= 32'd1073741827;
    else if (wr_en_i) rd_data_o <= wr_data_i;
  assign rd_error_o = 1'h0;
  assign rd_error_o_t0 = 1'h0;
endmodule

module paramoda05994007059a055454376e4d0aa9b8192775615auxy_prim_fifo_sync (clk_i, rst_ni, clr_i, wvalid_i, wready_o, wdata_i, rvalid_o, rready_i, rdata_o, full_o, depth_o, rready_i_t0, rvalid_o_t0, wdata_i_t0, wready_o_t0, wvalid_i_t0, clr_i_t0, depth_o_t0, full_o_t0, rdata_o_t0);
  wire [1:0] _000_;
  wire [1:0] _001_;
  wire [1:0] _002_;
  wire [1:0] _003_;
  wire _004_;
  wire _005_;
  wire _006_;
  wire _007_;
  wire [1:0] _008_;
  wire [1:0] _009_;
  wire [1:0] _010_;
  wire [1:0] _011_;
  wire _012_;
  wire _013_;
  wire _014_;
  wire _015_;
  wire _016_;
  wire _017_;
  wire _018_;
  wire _019_;
  wire _020_;
  wire _021_;
  wire [1:0] _022_;
  wire [1:0] _023_;
  wire _024_;
  wire _025_;
  wire _026_;
  wire [1:0] _027_;
  wire [1:0] _028_;
  wire _029_;
  wire [1:0] _030_;
  wire [1:0] _031_;
  wire [1:0] _032_;
  wire [1:0] _033_;
  wire [1:0] _034_;
  wire [1:0] _035_;
  wire _036_;
  wire _037_;
  wire _038_;
  wire _039_;
  wire [39:0] _040_;
  wire [39:0] _041_;
  wire _042_;
  wire _043_;
  wire _044_;
  wire _045_;
  wire _046_;
  wire _047_;
  wire _048_;
  wire _049_;
  wire _050_;
  wire [1:0] _051_;
  wire [1:0] _052_;
  wire _053_;
  wire _054_;
  wire _055_;
  wire _056_;
  wire _057_;
  wire _058_;
  wire _059_;
  wire _060_;
  wire _061_;
  wire _062_;
  wire _063_;
  wire _064_;
  wire _065_;
  wire _066_;
  wire _067_;
  wire _068_;
  wire _069_;
  wire _070_;
  wire _071_;
  wire _072_;
  wire _073_;
  wire [1:0] _074_;
  wire [1:0] _075_;
  wire [1:0] _076_;
  wire [39:0] _077_;
  wire [39:0] _078_;
  wire [39:0] _079_;
  wire [1:0] _080_;
  wire [1:0] _081_;
  wire [1:0] _082_;
  wire [1:0] _083_;
  wire [1:0] _084_;
  wire _085_;
  wire _086_;
  wire [1:0] _087_;
  wire [1:0] _088_;
  wire [1:0] _089_;
  wire _090_;
  wire [1:0] _091_;
  wire [1:0] _092_;
  wire [1:0] _093_;
  wire [1:0] _094_;
  wire [1:0] _095_;
  wire [1:0] _096_;
  wire [1:0] _097_;
  wire [1:0] _098_;
  wire [1:0] _099_;
  wire [1:0] _100_;
  wire [1:0] _101_;
  wire [1:0] _102_;
  wire [1:0] _103_;
  wire [1:0] _104_;
  wire [1:0] _105_;
  wire [1:0] _106_;
  wire [1:0] _107_;
  wire _108_;
  wire _109_;
  wire _110_;
  wire _111_;
  wire _112_;
  wire _113_;
  wire _114_;
  wire _115_;
  wire [39:0] _116_;
  wire [39:0] _117_;
  wire [39:0] _118_;
  wire [39:0] _119_;
  wire [39:0] _120_;
  wire [39:0] _121_;
  wire _122_;
  wire _123_;
  wire _124_;
  wire [1:0] _125_;
  wire [1:0] _126_;
  wire _127_;
  wire _128_;
  wire _129_;
  wire _130_;
  wire _131_;
  wire _132_;
  wire _133_;
  wire [1:0] _134_;
  wire [1:0] _135_;
  wire [1:0] _136_;
  wire [1:0] _137_;
  wire [39:0] _138_;
  wire [39:0] _139_;
  wire [39:0] _140_;
  wire [39:0] _141_;
  wire [1:0] _142_;
  wire [1:0] _143_;
  wire [1:0] _144_;
  wire [1:0] _145_;
  wire _146_;
  wire [1:0] _147_;
  wire _148_;
  wire [1:0] _149_;
  wire [1:0] _150_;
  wire [1:0] _151_;
  wire [1:0] _152_;
  wire [1:0] _153_;
  wire [1:0] _154_;
  wire [1:0] _155_;
  wire [1:0] _156_;
  wire [1:0] _157_;
  wire [1:0] _158_;
  wire [1:0] _159_;
  wire [1:0] _160_;
  wire [1:0] _161_;
  wire [1:0] _162_;
  wire [1:0] _163_;
  wire [1:0] _164_;
  wire _165_;
  wire _166_;
  wire _167_;
  wire _168_;
  wire _169_;
  wire _170_;
  wire _171_;
  wire _172_;
  wire [39:0] _173_;
  wire [39:0] _174_;
  wire [39:0] _175_;
  wire [39:0] _176_;
  wire [39:0] _177_;
  wire [39:0] _178_;
  wire _179_;
  wire [1:0] _180_;
  wire [1:0] _181_;
  wire [1:0] _182_;
  wire [39:0] _183_;
  wire [1:0] _184_;
  wire [1:0] _185_;
  wire [1:0] _186_;
  wire [1:0] _187_;
  wire [1:0] _188_;
  wire [1:0] _189_;
  wire [1:0] _190_;
  wire _191_;
  wire _192_;
  wire _193_;
  wire _194_;
  wire _195_;
  wire _196_;
  wire _197_;
  wire [1:0] _198_;
  wire [1:0] _199_;
  wire [1:0] _200_;
  wire [1:0] _201_;
  wire _202_;
  wire _203_;
  wire _204_;
  wire _205_;
  wire _206_;
  wire _207_;
  wire _208_;
  wire _209_;
  wire _210_;
  wire _211_;
  wire _212_;
  wire _213_;
  wire [1:0] _214_;
  wire [1:0] _215_;
  wire [1:0] _216_;
  wire [1:0] _217_;
  wire _218_;
  wire _219_;
  wire _220_;
  wire _221_;
  wire _222_;
  wire _223_;
  wire [1:0] _224_;
  input clk_i;
  wire clk_i;
  input clr_i;
  wire clr_i;
  input clr_i_t0;
  wire clr_i_t0;
  output depth_o;
  wire depth_o;
  output depth_o_t0;
  wire depth_o_t0;
  output full_o;
  wire full_o;
  output full_o_t0;
  wire full_o_t0;
  wire \gen_normal_fifo.empty ;
  wire \gen_normal_fifo.empty_t0 ;
  wire \gen_normal_fifo.fifo_empty ;
  wire \gen_normal_fifo.fifo_empty_t0 ;
  wire \gen_normal_fifo.fifo_incr_rptr ;
  wire \gen_normal_fifo.fifo_incr_rptr_t0 ;
  wire \gen_normal_fifo.fifo_incr_wptr ;
  wire \gen_normal_fifo.fifo_incr_wptr_t0 ;
  reg [1:0] \gen_normal_fifo.fifo_rptr ;
  reg [1:0] \gen_normal_fifo.fifo_rptr_t0 ;
  reg [1:0] \gen_normal_fifo.fifo_wptr ;
  reg [1:0] \gen_normal_fifo.fifo_wptr_t0 ;
  wire [39:0] \gen_normal_fifo.rdata_int ;
  wire [39:0] \gen_normal_fifo.rdata_int_t0 ;
  reg [39:0] \gen_normal_fifo.storage ;
  reg [39:0] \gen_normal_fifo.storage_t0 ;
  reg \gen_normal_fifo.under_rst ;
  reg \gen_normal_fifo.under_rst_t0 ;
  output [39:0] rdata_o;
  wire [39:0] rdata_o;
  output [39:0] rdata_o_t0;
  wire [39:0] rdata_o_t0;
  input rready_i;
  wire rready_i;
  input rready_i_t0;
  wire rready_i_t0;
  input rst_ni;
  wire rst_ni;
  output rvalid_o;
  wire rvalid_o;
  output rvalid_o_t0;
  wire rvalid_o_t0;
  input [39:0] wdata_i;
  wire [39:0] wdata_i;
  input [39:0] wdata_i_t0;
  wire [39:0] wdata_i_t0;
  output wready_o;
  wire wready_o;
  output wready_o_t0;
  wire wready_o_t0;
  input wvalid_i;
  wire wvalid_i;
  input wvalid_i_t0;
  wire wvalid_i_t0;
  assign _006_ = _220_ + \gen_normal_fifo.fifo_wptr [0];
  assign _008_ = \gen_normal_fifo.fifo_wptr  + 2'h1;
  assign _010_ = \gen_normal_fifo.fifo_rptr  + 2'h1;
  assign _012_ = wvalid_i & wready_o;
  assign \gen_normal_fifo.fifo_incr_wptr  = _012_ & _036_;
  assign _014_ = rvalid_o & rready_i;
  assign \gen_normal_fifo.fifo_incr_rptr  = _014_ & _036_;
  assign wready_o = _039_ & _036_;
  assign rvalid_o = _210_ & _036_;
  assign \gen_normal_fifo.empty  = \gen_normal_fifo.fifo_empty  & _213_;
  assign _020_ = ~ _221_;
  assign _022_ = ~ \gen_normal_fifo.fifo_wptr_t0 ;
  assign _023_ = ~ \gen_normal_fifo.fifo_rptr_t0 ;
  assign _049_ = _220_ & _020_;
  assign _051_ = \gen_normal_fifo.fifo_wptr  & _022_;
  assign _052_ = \gen_normal_fifo.fifo_rptr  & _023_;
  assign _196_ = _049_ + _050_;
  assign _198_ = _051_ + 2'h1;
  assign _200_ = _052_ + 2'h1;
  assign _122_ = _220_ | _221_;
  assign _125_ = \gen_normal_fifo.fifo_wptr  | \gen_normal_fifo.fifo_wptr_t0 ;
  assign _126_ = \gen_normal_fifo.fifo_rptr  | \gen_normal_fifo.fifo_rptr_t0 ;
  assign _197_ = _122_ + _123_;
  assign _199_ = _125_ + 2'h1;
  assign _201_ = _126_ + 2'h1;
  assign _179_ = _196_ ^ _197_;
  assign _180_ = _198_ ^ _199_;
  assign _181_ = _200_ ^ _201_;
  assign _124_ = _179_ | _221_;
  assign _009_ = _180_ | \gen_normal_fifo.fifo_wptr_t0 ;
  assign _011_ = _181_ | \gen_normal_fifo.fifo_rptr_t0 ;
  assign _007_ = _124_ | \gen_normal_fifo.fifo_wptr_t0 [0];
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) \gen_normal_fifo.under_rst_t0  <= 1'h0;
    else \gen_normal_fifo.under_rst_t0  <= _005_;
  assign _024_ = ~ _016_;
  assign _026_ = ~ _018_;
  assign _182_ = _002_ ^ \gen_normal_fifo.fifo_wptr ;
  assign _184_ = _000_ ^ \gen_normal_fifo.fifo_rptr ;
  assign _134_ = _003_ | \gen_normal_fifo.fifo_wptr_t0 ;
  assign _142_ = _001_ | \gen_normal_fifo.fifo_rptr_t0 ;
  assign _135_ = _182_ | _134_;
  assign _143_ = _184_ | _142_;
  assign _074_ = { _016_, _016_ } & _003_;
  assign _080_ = { _018_, _018_ } & _001_;
  assign _075_ = { _024_, _024_ } & \gen_normal_fifo.fifo_wptr_t0 ;
  assign _081_ = { _026_, _026_ } & \gen_normal_fifo.fifo_rptr_t0 ;
  assign _076_ = _135_ & { _017_, _017_ };
  assign _082_ = _143_ & { _019_, _019_ };
  assign _136_ = _074_ | _075_;
  assign _144_ = _080_ | _081_;
  assign _137_ = _136_ | _076_;
  assign _145_ = _144_ | _082_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) \gen_normal_fifo.fifo_wptr_t0  <= 2'h0;
    else \gen_normal_fifo.fifo_wptr_t0  <= _137_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) \gen_normal_fifo.fifo_rptr_t0  <= 2'h0;
    else \gen_normal_fifo.fifo_rptr_t0  <= _145_;
  assign _053_ = wvalid_i_t0 & wready_o;
  assign _056_ = _013_ & _036_;
  assign _059_ = rvalid_o_t0 & rready_i;
  assign _062_ = _015_ & _036_;
  assign _065_ = full_o_t0 & _036_;
  assign _068_ = \gen_normal_fifo.empty_t0  & _036_;
  assign _071_ = \gen_normal_fifo.fifo_empty_t0  & _213_;
  assign _054_ = wready_o_t0 & wvalid_i;
  assign _057_ = \gen_normal_fifo.under_rst_t0  & _012_;
  assign _060_ = rready_i_t0 & rvalid_o;
  assign _063_ = \gen_normal_fifo.under_rst_t0  & _014_;
  assign _066_ = \gen_normal_fifo.under_rst_t0  & _039_;
  assign _069_ = \gen_normal_fifo.under_rst_t0  & _210_;
  assign _055_ = wvalid_i_t0 & wready_o_t0;
  assign _058_ = _013_ & \gen_normal_fifo.under_rst_t0 ;
  assign _061_ = rvalid_o_t0 & rready_i_t0;
  assign _064_ = _015_ & \gen_normal_fifo.under_rst_t0 ;
  assign _067_ = full_o_t0 & \gen_normal_fifo.under_rst_t0 ;
  assign _070_ = \gen_normal_fifo.empty_t0  & \gen_normal_fifo.under_rst_t0 ;
  assign _127_ = _053_ | _054_;
  assign _128_ = _056_ | _057_;
  assign _129_ = _059_ | _060_;
  assign _130_ = _062_ | _063_;
  assign _131_ = _065_ | _066_;
  assign _132_ = _068_ | _069_;
  assign _133_ = _071_ | _072_;
  assign _013_ = _127_ | _055_;
  assign \gen_normal_fifo.fifo_incr_wptr_t0  = _128_ | _058_;
  assign _015_ = _129_ | _061_;
  assign \gen_normal_fifo.fifo_incr_rptr_t0  = _130_ | _064_;
  assign wready_o_t0 = _131_ | _067_;
  assign rvalid_o_t0 = _132_ | _070_;
  assign \gen_normal_fifo.empty_t0  = _133_ | _073_;
  assign _025_ = ~ \gen_normal_fifo.fifo_incr_wptr ;
  assign _138_ = wdata_i_t0 | \gen_normal_fifo.storage_t0 ;
  assign _139_ = _183_ | _138_;
  assign _077_ = { \gen_normal_fifo.fifo_incr_wptr , \gen_normal_fifo.fifo_incr_wptr , \gen_normal_fifo.fifo_incr_wptr , \gen_normal_fifo.fifo_incr_wptr , \gen_normal_fifo.fifo_incr_wptr , \gen_normal_fifo.fifo_incr_wptr , \gen_normal_fifo.fifo_incr_wptr , \gen_normal_fifo.fifo_incr_wptr , \gen_normal_fifo.fifo_incr_wptr , \gen_normal_fifo.fifo_incr_wptr , \gen_normal_fifo.fifo_incr_wptr , \gen_normal_fifo.fifo_incr_wptr , \gen_normal_fifo.fifo_incr_wptr , \gen_normal_fifo.fifo_incr_wptr , \gen_normal_fifo.fifo_incr_wptr , \gen_normal_fifo.fifo_incr_wptr , \gen_normal_fifo.fifo_incr_wptr , \gen_normal_fifo.fifo_incr_wptr , \gen_normal_fifo.fifo_incr_wptr , \gen_normal_fifo.fifo_incr_wptr , \gen_normal_fifo.fifo_incr_wptr , \gen_normal_fifo.fifo_incr_wptr , \gen_normal_fifo.fifo_incr_wptr , \gen_normal_fifo.fifo_incr_wptr , \gen_normal_fifo.fifo_incr_wptr , \gen_normal_fifo.fifo_incr_wptr , \gen_normal_fifo.fifo_incr_wptr , \gen_normal_fifo.fifo_incr_wptr , \gen_normal_fifo.fifo_incr_wptr , \gen_normal_fifo.fifo_incr_wptr , \gen_normal_fifo.fifo_incr_wptr , \gen_normal_fifo.fifo_incr_wptr , \gen_normal_fifo.fifo_incr_wptr , \gen_normal_fifo.fifo_incr_wptr , \gen_normal_fifo.fifo_incr_wptr , \gen_normal_fifo.fifo_incr_wptr , \gen_normal_fifo.fifo_incr_wptr , \gen_normal_fifo.fifo_incr_wptr , \gen_normal_fifo.fifo_incr_wptr , \gen_normal_fifo.fifo_incr_wptr  } & wdata_i_t0;
  assign _078_ = { _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_ } & \gen_normal_fifo.storage_t0 ;
  assign _079_ = _139_ & \gen_normal_fifo.fifo_incr_wptr_t0 ;
  assign _140_ = _077_ | _078_;
  assign _141_ = _140_ | _079_;
  always_ff @(posedge clk_i)
    \gen_normal_fifo.storage_t0  <= _141_;
  assign _045_ = | { \gen_normal_fifo.fifo_rptr_t0 [1], \gen_normal_fifo.fifo_wptr_t0 [1] };
  assign _046_ = | { \gen_normal_fifo.fifo_rptr_t0 , \gen_normal_fifo.fifo_wptr_t0  };
  assign _146_ = \gen_normal_fifo.fifo_wptr_t0 [1] | \gen_normal_fifo.fifo_rptr_t0 [1];
  assign _147_ = \gen_normal_fifo.fifo_wptr_t0  | \gen_normal_fifo.fifo_rptr_t0 ;
  assign _029_ = ~ _146_;
  assign _030_ = ~ _147_;
  assign _085_ = \gen_normal_fifo.fifo_wptr [1] & _029_;
  assign _087_ = \gen_normal_fifo.fifo_wptr  & _030_;
  assign _086_ = \gen_normal_fifo.fifo_rptr [1] & _029_;
  assign _088_ = _224_ & _030_;
  assign _089_ = \gen_normal_fifo.fifo_rptr  & _030_;
  assign _193_ = _085_ == _086_;
  assign _194_ = _087_ == _088_;
  assign _195_ = _087_ == _089_;
  assign _207_ = _193_ & _045_;
  assign full_o_t0 = _194_ & _046_;
  assign \gen_normal_fifo.fifo_empty_t0  = _195_ & _046_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) \gen_normal_fifo.fifo_wptr  <= 2'h0;
    else if (_016_) \gen_normal_fifo.fifo_wptr  <= _002_;
  always_ff @(posedge clk_i)
    if (\gen_normal_fifo.fifo_incr_wptr ) \gen_normal_fifo.storage  <= wdata_i;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) \gen_normal_fifo.fifo_rptr  <= 2'h0;
    else if (_018_) \gen_normal_fifo.fifo_rptr  <= _000_;
  assign _090_ = \gen_normal_fifo.fifo_empty_t0  & wvalid_i;
  assign _072_ = wvalid_i_t0 & \gen_normal_fifo.fifo_empty ;
  assign _073_ = \gen_normal_fifo.fifo_empty_t0  & wvalid_i_t0;
  assign _148_ = _090_ | _072_;
  assign _209_ = _148_ | _073_;
  assign _043_ = | { \gen_normal_fifo.fifo_incr_wptr_t0 , clr_i_t0 };
  assign _044_ = | { \gen_normal_fifo.fifo_incr_rptr_t0 , clr_i_t0 };
  assign _027_ = ~ { \gen_normal_fifo.fifo_incr_wptr_t0 , clr_i_t0 };
  assign _028_ = ~ { \gen_normal_fifo.fifo_incr_rptr_t0 , clr_i_t0 };
  assign _083_ = { \gen_normal_fifo.fifo_incr_wptr , clr_i } & _027_;
  assign _084_ = { \gen_normal_fifo.fifo_incr_rptr , clr_i } & _028_;
  assign _047_ = ! _083_;
  assign _048_ = ! _084_;
  assign _017_ = _047_ & _043_;
  assign _019_ = _048_ & _044_;
  assign _031_ = ~ { \gen_normal_fifo.fifo_rptr [0], \gen_normal_fifo.fifo_rptr [0] };
  assign _032_ = ~ { \gen_normal_fifo.fifo_incr_rptr , \gen_normal_fifo.fifo_incr_rptr  };
  assign _034_ = ~ { \gen_normal_fifo.fifo_wptr [0], \gen_normal_fifo.fifo_wptr [0] };
  assign _035_ = ~ { \gen_normal_fifo.fifo_incr_wptr , \gen_normal_fifo.fifo_incr_wptr  };
  assign _033_ = ~ { clr_i, clr_i };
  assign _036_ = ~ \gen_normal_fifo.under_rst ;
  assign _038_ = ~ _206_;
  assign _039_ = ~ full_o;
  assign _040_ = ~ { _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_ };
  assign _041_ = ~ { \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty  };
  assign _149_ = { \gen_normal_fifo.fifo_rptr_t0 [0], \gen_normal_fifo.fifo_rptr_t0 [0] } | _031_;
  assign _152_ = { \gen_normal_fifo.fifo_incr_rptr_t0 , \gen_normal_fifo.fifo_incr_rptr_t0  } | _032_;
  assign _158_ = { \gen_normal_fifo.fifo_wptr_t0 [0], \gen_normal_fifo.fifo_wptr_t0 [0] } | _034_;
  assign _161_ = { \gen_normal_fifo.fifo_incr_wptr_t0 , \gen_normal_fifo.fifo_incr_wptr_t0  } | _035_;
  assign _155_ = { clr_i_t0, clr_i_t0 } | _033_;
  assign _169_ = _207_ | _038_;
  assign _172_ = full_o_t0 | _039_;
  assign _173_ = { _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_ } | _040_;
  assign _176_ = { \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0  } | _041_;
  assign _150_ = { \gen_normal_fifo.fifo_rptr_t0 [0], \gen_normal_fifo.fifo_rptr_t0 [0] } | { \gen_normal_fifo.fifo_rptr [0], \gen_normal_fifo.fifo_rptr [0] };
  assign _153_ = { \gen_normal_fifo.fifo_incr_rptr_t0 , \gen_normal_fifo.fifo_incr_rptr_t0  } | { \gen_normal_fifo.fifo_incr_rptr , \gen_normal_fifo.fifo_incr_rptr  };
  assign _159_ = { \gen_normal_fifo.fifo_wptr_t0 [0], \gen_normal_fifo.fifo_wptr_t0 [0] } | { \gen_normal_fifo.fifo_wptr [0], \gen_normal_fifo.fifo_wptr [0] };
  assign _162_ = { \gen_normal_fifo.fifo_incr_wptr_t0 , \gen_normal_fifo.fifo_incr_wptr_t0  } | { \gen_normal_fifo.fifo_incr_wptr , \gen_normal_fifo.fifo_incr_wptr  };
  assign _156_ = { clr_i_t0, clr_i_t0 } | { clr_i, clr_i };
  assign _165_ = \gen_normal_fifo.under_rst_t0  | \gen_normal_fifo.under_rst ;
  assign _170_ = _207_ | _206_;
  assign _174_ = { _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_ } | { _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_ };
  assign _177_ = { \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0  } | { \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty  };
  assign _091_ = { \gen_normal_fifo.fifo_rptr_t0 [1], 1'h0 } & _149_;
  assign _094_ = 2'h0 & _152_;
  assign _097_ = _215_ & _155_;
  assign _100_ = { \gen_normal_fifo.fifo_wptr_t0 [1], 1'h0 } & _158_;
  assign _103_ = 2'h0 & _161_;
  assign _106_ = _217_ & _155_;
  assign _111_ = _007_ & _169_;
  assign _114_ = _223_ & _172_;
  assign _116_ = \gen_normal_fifo.storage_t0  & _173_;
  assign _119_ = \gen_normal_fifo.rdata_int_t0  & _176_;
  assign _092_ = _011_ & _150_;
  assign _095_ = _214_ & _153_;
  assign _101_ = _009_ & _159_;
  assign _104_ = _216_ & _162_;
  assign _098_ = 2'h0 & _156_;
  assign _108_ = \gen_normal_fifo.under_rst_t0  & _165_;
  assign _112_ = _219_ & _170_;
  assign _117_ = wdata_i_t0 & _174_;
  assign _120_ = 40'h0000000000 & _177_;
  assign _151_ = _091_ | _092_;
  assign _154_ = _094_ | _095_;
  assign _157_ = _097_ | _098_;
  assign _160_ = _100_ | _101_;
  assign _163_ = _103_ | _104_;
  assign _164_ = _106_ | _098_;
  assign _171_ = _111_ | _112_;
  assign _175_ = _116_ | _117_;
  assign _178_ = _119_ | _120_;
  assign _185_ = { _212_, 1'h0 } ^ _010_;
  assign _188_ = { _211_, 1'h0 } ^ _008_;
  assign _192_ = _006_ ^ _218_;
  assign _183_ = \gen_normal_fifo.storage  ^ wdata_i;
  assign _093_ = { \gen_normal_fifo.fifo_rptr_t0 [0], \gen_normal_fifo.fifo_rptr_t0 [0] } & _185_;
  assign _096_ = { \gen_normal_fifo.fifo_incr_rptr_t0 , \gen_normal_fifo.fifo_incr_rptr_t0  } & _186_;
  assign _099_ = { clr_i_t0, clr_i_t0 } & _187_;
  assign _102_ = { \gen_normal_fifo.fifo_wptr_t0 [0], \gen_normal_fifo.fifo_wptr_t0 [0] } & _188_;
  assign _105_ = { \gen_normal_fifo.fifo_incr_wptr_t0 , \gen_normal_fifo.fifo_incr_wptr_t0  } & _189_;
  assign _107_ = { clr_i_t0, clr_i_t0 } & _190_;
  assign _109_ = \gen_normal_fifo.under_rst_t0  & _036_;
  assign _113_ = _207_ & _192_;
  assign _115_ = full_o_t0 & _042_;
  assign _118_ = { _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_ } & _183_;
  assign _121_ = { \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0  } & \gen_normal_fifo.rdata_int ;
  assign _214_ = _093_ | _151_;
  assign _215_ = _096_ | _154_;
  assign _001_ = _099_ | _157_;
  assign _216_ = _102_ | _160_;
  assign _217_ = _105_ | _163_;
  assign _003_ = _107_ | _164_;
  assign _005_ = _109_ | _108_;
  assign _223_ = _113_ | _171_;
  assign depth_o_t0 = _115_ | _114_;
  assign \gen_normal_fifo.rdata_int_t0  = _118_ | _175_;
  assign rdata_o_t0 = _121_ | _178_;
  assign _016_ = | { \gen_normal_fifo.fifo_incr_wptr , clr_i };
  assign _018_ = | { \gen_normal_fifo.fifo_incr_rptr , clr_i };
  assign _042_ = ~ _222_;
  assign _021_ = ~ \gen_normal_fifo.fifo_wptr_t0 [0];
  assign _037_ = ~ \gen_normal_fifo.fifo_rptr_t0 [0];
  assign _050_ = \gen_normal_fifo.fifo_wptr [0] & _021_;
  assign _110_ = \gen_normal_fifo.fifo_rptr [0] & _037_;
  assign _123_ = \gen_normal_fifo.fifo_wptr [0] | \gen_normal_fifo.fifo_wptr_t0 [0];
  assign _166_ = \gen_normal_fifo.fifo_rptr [0] | \gen_normal_fifo.fifo_rptr_t0 [0];
  assign _202_ = _123_ - _110_;
  assign _204_ = 1'h1 - _110_;
  assign _203_ = _050_ - _166_;
  assign _205_ = 1'h1 - _166_;
  assign _191_ = _202_ ^ _203_;
  assign _168_ = _204_ ^ _205_;
  assign _167_ = _191_ | \gen_normal_fifo.fifo_wptr_t0 [0];
  assign _219_ = _167_ | \gen_normal_fifo.fifo_rptr_t0 [0];
  assign _221_ = _168_ | \gen_normal_fifo.fifo_rptr_t0 [0];
  assign _206_ = \gen_normal_fifo.fifo_wptr [1] == \gen_normal_fifo.fifo_rptr [1];
  assign full_o = \gen_normal_fifo.fifo_wptr  == _224_;
  assign \gen_normal_fifo.fifo_empty  = \gen_normal_fifo.fifo_wptr  == \gen_normal_fifo.fifo_rptr ;
  assign _208_ = \gen_normal_fifo.fifo_empty  && wvalid_i;
  assign _210_ = ~ \gen_normal_fifo.empty ;
  assign _211_ = ~ \gen_normal_fifo.fifo_wptr [1];
  assign _212_ = ~ \gen_normal_fifo.fifo_rptr [1];
  assign _213_ = ~ wvalid_i;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) \gen_normal_fifo.under_rst  <= 1'h1;
    else \gen_normal_fifo.under_rst  <= _004_;
  assign _186_ = \gen_normal_fifo.fifo_rptr [0] ? _010_ : { _212_, 1'h0 };
  assign _187_ = \gen_normal_fifo.fifo_incr_rptr  ? _186_ : 2'hx;
  assign _000_ = clr_i ? 2'h0 : _187_;
  assign _189_ = \gen_normal_fifo.fifo_wptr [0] ? _008_ : { _211_, 1'h0 };
  assign _190_ = \gen_normal_fifo.fifo_incr_wptr  ? _189_ : 2'hx;
  assign _002_ = clr_i ? 2'h0 : _190_;
  assign _004_ = \gen_normal_fifo.under_rst  ? _036_ : 1'h0;
  assign _218_ = \gen_normal_fifo.fifo_wptr [0] - \gen_normal_fifo.fifo_rptr [0];
  assign _220_ = 1'h1 - \gen_normal_fifo.fifo_rptr [0];
  assign _222_ = _206_ ? _218_ : _006_;
  assign depth_o = full_o ? 1'h1 : _222_;
  assign \gen_normal_fifo.rdata_int  = _208_ ? wdata_i : \gen_normal_fifo.storage ;
  assign rdata_o = \gen_normal_fifo.empty  ? 40'h0000000000 : \gen_normal_fifo.rdata_int ;
  assign _224_ = \gen_normal_fifo.fifo_rptr  ^ 2'h2;
endmodule

module paramoda7b3f37e1f713a4d0901b62b3f601f61ae6218e0auxy_ibex_cs_registers (clk_i, rst_ni, hart_id_i, priv_mode_id_o, priv_mode_if_o, priv_mode_lsu_o, csr_mstatus_tw_o, csr_mtvec_o, csr_mtvec_init_i, boot_addr_i, csr_access_i, csr_addr_i, csr_wdata_i, csr_op_i, csr_op_en_i, csr_rdata_o, irq_software_i, irq_timer_i, irq_external_i, irq_fast_i, nmi_mode_i
, irq_pending_o, irqs_o, csr_mstatus_mie_o, csr_mepc_o, csr_pmp_cfg_o, csr_pmp_addr_o, csr_pmp_mseccfg_o, debug_mode_i, debug_cause_i, debug_csr_save_i, csr_depc_o, debug_single_step_o, debug_ebreakm_o, debug_ebreaku_o, trigger_match_o, pc_if_i, pc_id_i, pc_wb_i, data_ind_timing_o, dummy_instr_en_o, dummy_instr_mask_o
, dummy_instr_seed_en_o, dummy_instr_seed_o, icache_enable_o, csr_shadow_err_o, csr_save_if_i, csr_save_id_i, csr_save_wb_i, csr_restore_mret_i, csr_restore_dret_i, csr_save_cause_i, csr_mcause_i, csr_mtval_i, illegal_csr_insn_o, instr_ret_i, instr_ret_compressed_i, iside_wait_i, jump_i, branch_i, branch_taken_i, mem_load_i, mem_store_i
, dside_wait_i, mul_wait_i, div_wait_i, boot_addr_i_t0, branch_i_t0, branch_taken_i_t0, pc_id_i_t0, csr_access_i_t0, csr_addr_i_t0, csr_depc_o_t0, csr_mcause_i_t0, csr_mepc_o_t0, csr_mstatus_mie_o_t0, csr_mstatus_tw_o_t0, csr_mtval_i_t0, csr_mtvec_init_i_t0, csr_mtvec_o_t0, csr_op_en_i_t0, csr_op_i_t0, csr_pmp_addr_o_t0, csr_pmp_cfg_o_t0
, csr_pmp_mseccfg_o_t0, csr_rdata_o_t0, csr_restore_dret_i_t0, csr_restore_mret_i_t0, csr_save_cause_i_t0, csr_save_id_i_t0, csr_save_if_i_t0, csr_save_wb_i_t0, csr_shadow_err_o_t0, csr_wdata_i_t0, data_ind_timing_o_t0, debug_cause_i_t0, debug_csr_save_i_t0, debug_ebreakm_o_t0, debug_ebreaku_o_t0, debug_mode_i_t0, debug_single_step_o_t0, div_wait_i_t0, dside_wait_i_t0, dummy_instr_en_o_t0, dummy_instr_mask_o_t0
, dummy_instr_seed_en_o_t0, dummy_instr_seed_o_t0, hart_id_i_t0, icache_enable_o_t0, illegal_csr_insn_o_t0, instr_ret_compressed_i_t0, instr_ret_i_t0, irq_external_i_t0, irq_fast_i_t0, irq_pending_o_t0, irq_software_i_t0, irq_timer_i_t0, irqs_o_t0, iside_wait_i_t0, jump_i_t0, mem_load_i_t0, mem_store_i_t0, mul_wait_i_t0, nmi_mode_i_t0, pc_if_i_t0, pc_wb_i_t0
, priv_mode_id_o_t0, priv_mode_if_o_t0, priv_mode_lsu_o_t0, trigger_match_o_t0);
  wire [31:0] _0000_;
  wire [31:0] _0001_;
  wire _0002_;
  wire _0003_;
  wire _0004_;
  wire _0005_;
  wire _0006_;
  wire _0007_;
  wire _0008_;
  wire _0009_;
  wire [5:0] _0010_;
  wire [5:0] _0011_;
  wire _0012_;
  wire _0013_;
  wire _0014_;
  wire _0015_;
  wire [63:0] _0016_;
  wire [63:0] _0017_;
  wire [31:0] _0018_;
  wire [31:0] _0019_;
  wire _0020_;
  wire _0021_;
  wire [31:0] _0022_;
  wire [31:0] _0023_;
  wire _0024_;
  wire _0025_;
  wire [31:0] _0026_;
  wire [31:0] _0027_;
  wire _0028_;
  wire _0029_;
  wire _0030_;
  wire _0031_;
  wire _0032_;
  wire _0033_;
  wire [31:0] _0034_;
  wire [31:0] _0035_;
  wire [5:0] _0036_;
  wire [5:0] _0037_;
  wire _0038_;
  wire _0039_;
  wire _0040_;
  wire _0041_;
  wire [31:0] _0042_;
  wire [31:0] _0043_;
  wire _0044_;
  wire _0045_;
  wire [31:0] _0046_;
  wire [31:0] _0047_;
  wire [31:0] _0048_;
  wire [31:0] _0049_;
  wire _0050_;
  wire _0051_;
  wire _0052_;
  wire _0053_;
  wire _0054_;
  wire _0055_;
  wire [5:0] _0056_;
  wire [5:0] _0057_;
  wire _0058_;
  wire _0059_;
  wire [31:0] _0060_;
  wire [31:0] _0061_;
  wire _0062_;
  wire _0063_;
  wire _0064_;
  wire _0065_;
  wire [1:0] _0066_;
  wire [1:0] _0067_;
  wire [5:0] _0068_;
  wire [5:0] _0069_;
  wire [31:0] _0070_;
  wire [31:0] _0071_;
  wire _0072_;
  wire [1:0] _0073_;
  wire [1:0] _0074_;
  wire [31:0] _0075_;
  wire [31:0] _0076_;
  wire _0077_;
  wire _0078_;
  wire _0079_;
  wire _0080_;
  wire [5:0] _0081_;
  wire [5:0] _0082_;
  wire _0083_;
  wire _0084_;
  wire [31:0] _0085_;
  wire [31:0] _0086_;
  wire _0087_;
  wire _0088_;
  wire _0089_;
  wire _0090_;
  wire _0091_;
  wire _0092_;
  wire _0093_;
  wire _0094_;
  wire _0095_;
  wire _0096_;
  wire [3:0] _0097_;
  wire [3:0] _0098_;
  wire _0099_;
  wire _0100_;
  wire _0101_;
  wire _0102_;
  wire [1:0] _0103_;
  wire [1:0] _0104_;
  wire _0105_;
  wire _0106_;
  wire _0107_;
  wire _0108_;
  wire [3:0] _0109_;
  wire [3:0] _0110_;
  wire [2:0] _0111_;
  wire [2:0] _0112_;
  wire [2:0] _0113_;
  wire [2:0] _0114_;
  wire [31:0] _0115_;
  wire [31:0] _0116_;
  wire [31:0] _0117_;
  wire [31:0] _0118_;
  wire _0119_;
  wire _0120_;
  wire _0121_;
  wire _0122_;
  wire _0123_;
  wire _0124_;
  wire _0125_;
  wire _0126_;
  wire _0127_;
  wire _0128_;
  wire _0129_;
  wire _0130_;
  wire _0131_;
  wire _0132_;
  wire _0133_;
  wire _0134_;
  wire _0135_;
  wire _0136_;
  wire _0137_;
  wire _0138_;
  wire _0139_;
  wire _0140_;
  wire _0141_;
  wire _0142_;
  wire _0143_;
  wire _0144_;
  wire _0145_;
  wire _0146_;
  wire _0147_;
  wire _0148_;
  wire _0149_;
  wire _0150_;
  wire _0151_;
  wire _0152_;
  wire _0153_;
  wire _0154_;
  wire _0155_;
  wire _0156_;
  wire _0157_;
  wire _0158_;
  wire _0159_;
  wire _0160_;
  wire _0161_;
  wire _0162_;
  wire _0163_;
  wire _0164_;
  wire [130:0] _0165_;
  wire [3:0] _0166_;
  wire [19:0] _0167_;
  wire [1:0] _0168_;
  wire [1:0] _0169_;
  wire _0170_;
  wire _0171_;
  wire _0172_;
  wire _0173_;
  wire _0174_;
  wire _0175_;
  wire _0176_;
  wire _0177_;
  wire _0178_;
  wire _0179_;
  wire _0180_;
  wire _0181_;
  wire _0182_;
  wire _0183_;
  wire _0184_;
  wire _0185_;
  wire _0186_;
  wire _0187_;
  wire _0188_;
  wire _0189_;
  wire [2:0] _0190_;
  wire [2:0] _0191_;
  wire [32:0] _0192_;
  wire [2:0] _0193_;
  wire [36:0] _0194_;
  wire [63:0] _0195_;
  wire [2:0] _0196_;
  wire [3:0] _0197_;
  wire [67:0] _0198_;
  wire [21:0] _0199_;
  wire [2:0] _0200_;
  wire [24:0] _0201_;
  wire [62:0] _0202_;
  wire [3:0] _0203_;
  wire [66:0] _0204_;
  wire [62:0] _0205_;
  wire [65:0] _0206_;
  wire [64:0] _0207_;
  wire [2:0] _0208_;
  wire [63:0] _0209_;
  wire [60:0] _0210_;
  wire [2:0] _0211_;
  wire [33:0] _0212_;
  wire [3:0] _0213_;
  wire [37:0] _0214_;
  wire [62:0] _0215_;
  wire [2:0] _0216_;
  wire [65:0] _0217_;
  wire [31:0] _0218_;
  wire [31:0] _0219_;
  wire _0220_;
  wire _0221_;
  wire _0222_;
  wire _0223_;
  wire _0224_;
  wire _0225_;
  wire _0226_;
  wire _0227_;
  wire _0228_;
  wire [2:0] _0229_;
  wire [2:0] _0230_;
  wire [2:0] _0231_;
  wire [2:0] _0232_;
  wire [2:0] _0233_;
  wire [2:0] _0234_;
  wire [2:0] _0235_;
  wire [2:0] _0236_;
  wire [2:0] _0237_;
  wire [2:0] _0238_;
  wire [2:0] _0239_;
  wire [2:0] _0240_;
  wire [2:0] _0241_;
  wire [2:0] _0242_;
  wire [2:0] _0243_;
  wire _0244_;
  wire _0245_;
  wire _0246_;
  wire _0247_;
  wire _0248_;
  wire [2:0] _0249_;
  wire [2:0] _0250_;
  wire [2:0] _0251_;
  wire [2:0] _0252_;
  wire [2:0] _0253_;
  wire [2:0] _0254_;
  wire [2:0] _0255_;
  wire [2:0] _0256_;
  wire [2:0] _0257_;
  wire [2:0] _0258_;
  wire [2:0] _0259_;
  wire [2:0] _0260_;
  wire [31:0] _0261_;
  wire [31:0] _0262_;
  wire [31:0] _0263_;
  wire [31:0] _0264_;
  wire [31:0] _0265_;
  wire [31:0] _0266_;
  wire [31:0] _0267_;
  wire [31:0] _0268_;
  wire [31:0] _0269_;
  wire [31:0] _0270_;
  wire [31:0] _0271_;
  wire [31:0] _0272_;
  wire _0273_;
  wire _0274_;
  wire _0275_;
  wire _0276_;
  wire _0277_;
  wire _0278_;
  wire _0279_;
  wire [63:0] _0280_;
  wire [63:0] _0281_;
  wire [63:0] _0282_;
  wire [63:0] _0283_;
  wire [63:0] _0284_;
  wire [63:0] _0285_;
  wire [63:0] _0286_;
  wire [63:0] _0287_;
  wire [63:0] _0288_;
  wire [63:0] _0289_;
  wire [63:0] _0290_;
  wire [63:0] _0291_;
  wire [8:0] _0292_;
  wire [8:0] _0293_;
  wire [8:0] _0294_;
  wire [8:0] _0295_;
  wire [8:0] _0296_;
  wire [8:0] _0297_;
  wire [8:0] _0298_;
  wire [8:0] _0299_;
  wire [8:0] _0300_;
  wire [8:0] _0301_;
  wire [8:0] _0302_;
  wire [8:0] _0303_;
  wire [8:0] _0304_;
  wire [8:0] _0305_;
  wire [8:0] _0306_;
  wire [8:0] _0307_;
  wire [8:0] _0308_;
  wire [8:0] _0309_;
  wire [2:0] _0310_;
  wire [2:0] _0311_;
  wire [2:0] _0312_;
  wire [2:0] _0313_;
  wire [2:0] _0314_;
  wire [2:0] _0315_;
  wire [2:0] _0316_;
  wire [2:0] _0317_;
  wire [2:0] _0318_;
  wire [2:0] _0319_;
  wire [2:0] _0320_;
  wire [2:0] _0321_;
  wire [2:0] _0322_;
  wire [2:0] _0323_;
  wire _0324_;
  wire [2:0] _0325_;
  wire [2:0] _0326_;
  wire [2:0] _0327_;
  wire [2:0] _0328_;
  wire [2:0] _0329_;
  wire _0330_;
  wire _0331_;
  wire _0332_;
  wire _0333_;
  wire _0334_;
  wire _0335_;
  wire [1:0] _0336_;
  wire [31:0] _0337_;
  wire _0338_;
  wire _0339_;
  wire _0340_;
  wire _0341_;
  wire [30:0] _0342_;
  wire _0343_;
  wire [1:0] _0344_;
  wire [1:0] _0345_;
  wire [31:0] _0346_;
  wire [31:0] _0347_;
  wire [31:0] _0348_;
  wire _0349_;
  wire _0350_;
  wire _0351_;
  wire _0352_;
  wire [31:0] _0353_;
  wire [31:0] _0354_;
  wire _0355_;
  wire _0356_;
  wire _0357_;
  wire _0358_;
  wire [1:0] _0359_;
  wire _0360_;
  wire _0361_;
  wire _0362_;
  wire _0363_;
  wire [31:0] _0364_;
  wire [1:0] _0365_;
  wire [2:0] _0366_;
  wire [2:0] _0367_;
  wire [2:0] _0368_;
  wire [5:0] _0369_;
  wire [5:0] _0370_;
  wire _0371_;
  wire [31:0] _0372_;
  wire [1:0] _0373_;
  wire _0374_;
  wire [31:0] _0375_;
  wire [2:0] _0376_;
  wire [1:0] _0377_;
  wire [5:0] _0378_;
  wire [3:0] _0379_;
  wire [31:0] _0380_;
  wire [31:0] _0381_;
  wire [31:0] _0382_;
  wire [31:0] _0383_;
  wire [1:0] _0384_;
  wire [5:0] _0385_;
  wire [5:0] _0386_;
  wire [5:0] _0387_;
  wire [31:0] _0388_;
  wire [31:0] _0389_;
  wire [1:0] _0390_;
  wire [1:0] _0391_;
  wire [3:0] _0392_;
  wire [1:0] _0393_;
  wire [11:0] _0394_;
  wire [1:0] _0395_;
  wire [1:0] _0396_;
  wire [1:0] _0397_;
  wire [31:0] _0398_;
  wire [31:0] _0399_;
  wire _0400_;
  wire [31:0] _0401_;
  wire [5:0] _0402_;
  wire [30:0] _0403_;
  wire [28:0] _0404_;
  wire [11:0] _0405_;
  wire [4:0] _0406_;
  wire [30:0] _0407_;
  wire [2:0] _0408_;
  wire [17:0] _0409_;
  wire [31:0] _0410_;
  wire [1:0] _0411_;
  wire _0412_;
  wire _0413_;
  wire _0414_;
  wire _0415_;
  wire _0416_;
  wire _0417_;
  wire _0418_;
  wire _0419_;
  wire _0420_;
  wire _0421_;
  wire _0422_;
  wire _0423_;
  wire _0424_;
  wire _0425_;
  wire [31:0] _0426_;
  wire [31:0] _0427_;
  wire _0428_;
  wire _0429_;
  wire _0430_;
  wire _0431_;
  wire _0432_;
  wire _0433_;
  wire _0434_;
  wire _0435_;
  wire _0436_;
  wire _0437_;
  wire _0438_;
  wire _0439_;
  wire _0440_;
  wire _0441_;
  wire _0442_;
  wire _0443_;
  wire _0444_;
  wire _0445_;
  wire _0446_;
  wire _0447_;
  wire _0448_;
  wire _0449_;
  wire _0450_;
  wire _0451_;
  wire _0452_;
  wire _0453_;
  wire _0454_;
  wire _0455_;
  wire _0456_;
  wire _0457_;
  wire _0458_;
  wire _0459_;
  wire _0460_;
  wire _0461_;
  wire _0462_;
  wire _0463_;
  wire _0464_;
  wire _0465_;
  wire _0466_;
  wire _0467_;
  wire _0468_;
  wire _0469_;
  wire _0470_;
  wire _0471_;
  wire _0472_;
  wire _0473_;
  wire _0474_;
  wire _0475_;
  wire _0476_;
  wire _0477_;
  wire _0478_;
  wire _0479_;
  wire _0480_;
  wire _0481_;
  wire _0482_;
  wire _0483_;
  wire _0484_;
  wire _0485_;
  wire _0486_;
  wire _0487_;
  wire _0488_;
  wire _0489_;
  wire _0490_;
  wire _0491_;
  wire _0492_;
  wire _0493_;
  wire _0494_;
  wire _0495_;
  wire _0496_;
  wire _0497_;
  wire _0498_;
  wire _0499_;
  wire _0500_;
  wire _0501_;
  wire _0502_;
  wire _0503_;
  wire _0504_;
  wire _0505_;
  wire _0506_;
  wire _0507_;
  wire _0508_;
  wire _0509_;
  wire _0510_;
  wire _0511_;
  wire _0512_;
  wire _0513_;
  wire _0514_;
  wire _0515_;
  wire _0516_;
  wire _0517_;
  wire _0518_;
  wire _0519_;
  wire _0520_;
  wire _0521_;
  wire _0522_;
  wire _0523_;
  wire _0524_;
  wire _0525_;
  wire _0526_;
  wire _0527_;
  wire _0528_;
  wire _0529_;
  wire _0530_;
  wire _0531_;
  wire _0532_;
  wire _0533_;
  wire _0534_;
  wire _0535_;
  wire _0536_;
  wire _0537_;
  wire _0538_;
  wire _0539_;
  wire _0540_;
  wire _0541_;
  wire _0542_;
  wire _0543_;
  wire _0544_;
  wire _0545_;
  wire _0546_;
  wire _0547_;
  wire _0548_;
  wire _0549_;
  wire _0550_;
  wire _0551_;
  wire _0552_;
  wire _0553_;
  wire _0554_;
  wire _0555_;
  wire _0556_;
  wire _0557_;
  wire _0558_;
  wire _0559_;
  wire _0560_;
  wire _0561_;
  wire _0562_;
  wire _0563_;
  wire _0564_;
  wire _0565_;
  wire _0566_;
  wire _0567_;
  wire _0568_;
  wire _0569_;
  wire _0570_;
  wire [31:0] _0571_;
  wire _0572_;
  wire _0573_;
  wire _0574_;
  wire [31:0] _0575_;
  wire [31:0] _0576_;
  wire [31:0] _0577_;
  wire _0578_;
  wire _0579_;
  wire _0580_;
  wire _0581_;
  wire _0582_;
  wire _0583_;
  wire [17:0] _0584_;
  wire [17:0] _0585_;
  wire [17:0] _0586_;
  wire _0587_;
  wire _0588_;
  wire _0589_;
  wire _0590_;
  wire _0591_;
  wire _0592_;
  wire _0593_;
  wire _0594_;
  wire _0595_;
  wire _0596_;
  wire _0597_;
  wire _0598_;
  wire _0599_;
  wire _0600_;
  wire _0601_;
  wire _0602_;
  wire _0603_;
  wire _0604_;
  wire _0605_;
  wire _0606_;
  wire _0607_;
  wire _0608_;
  wire _0609_;
  wire _0610_;
  wire _0611_;
  wire _0612_;
  wire _0613_;
  wire _0614_;
  wire _0615_;
  wire _0616_;
  wire _0617_;
  wire _0618_;
  wire _0619_;
  wire _0620_;
  wire _0621_;
  wire _0622_;
  wire _0623_;
  wire _0624_;
  wire _0625_;
  wire _0626_;
  wire _0627_;
  wire _0628_;
  wire _0629_;
  wire _0630_;
  wire _0631_;
  wire _0632_;
  wire _0633_;
  wire _0634_;
  wire _0635_;
  wire _0636_;
  wire _0637_;
  wire _0638_;
  wire _0639_;
  wire _0640_;
  wire [11:0] _0641_;
  wire [11:0] _0642_;
  wire [11:0] _0643_;
  wire [130:0] _0644_;
  wire [3:0] _0645_;
  wire [19:0] _0646_;
  wire [1:0] _0647_;
  wire [1:0] _0648_;
  wire _0649_;
  wire _0650_;
  wire _0651_;
  wire _0652_;
  wire _0653_;
  wire _0654_;
  wire _0655_;
  wire _0656_;
  wire _0657_;
  wire _0658_;
  wire _0659_;
  wire _0660_;
  wire _0661_;
  wire _0662_;
  wire _0663_;
  wire _0664_;
  wire _0665_;
  wire _0666_;
  wire _0667_;
  wire _0668_;
  wire _0669_;
  wire _0670_;
  wire _0671_;
  wire _0672_;
  wire _0673_;
  wire _0674_;
  wire _0675_;
  wire _0676_;
  wire _0677_;
  wire _0678_;
  wire _0679_;
  wire _0680_;
  wire _0681_;
  wire _0682_;
  wire _0683_;
  wire _0684_;
  wire _0685_;
  wire _0686_;
  wire _0687_;
  wire _0688_;
  wire _0689_;
  wire _0690_;
  wire _0691_;
  wire _0692_;
  wire _0693_;
  wire _0694_;
  wire _0695_;
  wire _0696_;
  wire [2:0] _0697_;
  wire [2:0] _0698_;
  wire [32:0] _0699_;
  wire [2:0] _0700_;
  wire [36:0] _0701_;
  wire [63:0] _0702_;
  wire [2:0] _0703_;
  wire [3:0] _0704_;
  wire [67:0] _0705_;
  wire [21:0] _0706_;
  wire [2:0] _0707_;
  wire [24:0] _0708_;
  wire [62:0] _0709_;
  wire [3:0] _0710_;
  wire [66:0] _0711_;
  wire [62:0] _0712_;
  wire [65:0] _0713_;
  wire [64:0] _0714_;
  wire [2:0] _0715_;
  wire [63:0] _0716_;
  wire [60:0] _0717_;
  wire [2:0] _0718_;
  wire [33:0] _0719_;
  wire [3:0] _0720_;
  wire [37:0] _0721_;
  wire [62:0] _0722_;
  wire [2:0] _0723_;
  wire [65:0] _0724_;
  wire [31:0] _0725_;
  wire [31:0] _0726_;
  wire [31:0] _0727_;
  wire [31:0] _0728_;
  wire [31:0] _0729_;
  wire [31:0] _0730_;
  wire _0731_;
  wire _0732_;
  wire _0733_;
  wire _0734_;
  wire _0735_;
  wire _0736_;
  wire _0737_;
  wire _0738_;
  wire _0739_;
  wire _0740_;
  wire _0741_;
  wire _0742_;
  wire _0743_;
  wire _0744_;
  wire _0745_;
  wire _0746_;
  wire _0747_;
  wire _0748_;
  wire _0749_;
  wire _0750_;
  wire _0751_;
  wire _0752_;
  wire _0753_;
  wire _0754_;
  wire _0755_;
  wire _0756_;
  wire _0757_;
  wire _0758_;
  wire _0759_;
  wire _0760_;
  wire _0761_;
  wire _0762_;
  wire _0763_;
  wire _0764_;
  wire _0765_;
  wire _0766_;
  wire _0767_;
  wire _0768_;
  wire _0769_;
  wire _0770_;
  wire _0771_;
  wire _0772_;
  wire _0773_;
  wire [2:0] _0774_;
  wire [2:0] _0775_;
  wire [2:0] _0776_;
  wire [2:0] _0777_;
  wire [2:0] _0778_;
  wire [2:0] _0779_;
  wire [2:0] _0780_;
  wire [2:0] _0781_;
  wire [2:0] _0782_;
  wire [2:0] _0783_;
  wire [2:0] _0784_;
  wire [2:0] _0785_;
  wire [2:0] _0786_;
  wire [2:0] _0787_;
  wire [2:0] _0788_;
  wire [2:0] _0789_;
  wire [2:0] _0790_;
  wire [2:0] _0791_;
  wire [2:0] _0792_;
  wire [2:0] _0793_;
  wire [2:0] _0794_;
  wire [2:0] _0795_;
  wire [2:0] _0796_;
  wire [2:0] _0797_;
  wire [2:0] _0798_;
  wire [2:0] _0799_;
  wire [2:0] _0800_;
  wire [2:0] _0801_;
  wire [2:0] _0802_;
  wire [2:0] _0803_;
  wire [2:0] _0804_;
  wire [2:0] _0805_;
  wire [2:0] _0806_;
  wire [2:0] _0807_;
  wire [2:0] _0808_;
  wire [2:0] _0809_;
  wire [2:0] _0810_;
  wire [2:0] _0811_;
  wire [2:0] _0812_;
  wire [2:0] _0813_;
  wire [2:0] _0814_;
  wire [2:0] _0815_;
  wire [2:0] _0816_;
  wire [2:0] _0817_;
  wire [2:0] _0818_;
  wire _0819_;
  wire _0820_;
  wire _0821_;
  wire _0822_;
  wire _0823_;
  wire _0824_;
  wire _0825_;
  wire _0826_;
  wire _0827_;
  wire _0828_;
  wire _0829_;
  wire _0830_;
  wire _0831_;
  wire _0832_;
  wire _0833_;
  wire _0834_;
  wire _0835_;
  wire _0836_;
  wire _0837_;
  wire _0838_;
  wire _0839_;
  wire _0840_;
  wire _0841_;
  wire _0842_;
  wire _0843_;
  wire _0844_;
  wire _0845_;
  wire _0846_;
  wire _0847_;
  wire _0848_;
  wire _0849_;
  wire _0850_;
  wire _0851_;
  wire _0852_;
  wire _0853_;
  wire _0854_;
  wire _0855_;
  wire _0856_;
  wire _0857_;
  wire _0858_;
  wire _0859_;
  wire _0860_;
  wire _0861_;
  wire _0862_;
  wire _0863_;
  wire _0864_;
  wire _0865_;
  wire _0866_;
  wire _0867_;
  wire _0868_;
  wire [2:0] _0869_;
  wire [2:0] _0870_;
  wire [2:0] _0871_;
  wire [2:0] _0872_;
  wire [2:0] _0873_;
  wire [2:0] _0874_;
  wire [2:0] _0875_;
  wire [2:0] _0876_;
  wire [2:0] _0877_;
  wire [2:0] _0878_;
  wire [2:0] _0879_;
  wire [2:0] _0880_;
  wire [2:0] _0881_;
  wire [2:0] _0882_;
  wire [2:0] _0883_;
  wire [2:0] _0884_;
  wire [2:0] _0885_;
  wire [2:0] _0886_;
  wire [2:0] _0887_;
  wire [2:0] _0888_;
  wire [2:0] _0889_;
  wire [2:0] _0890_;
  wire [2:0] _0891_;
  wire [2:0] _0892_;
  wire [2:0] _0893_;
  wire [2:0] _0894_;
  wire [2:0] _0895_;
  wire [2:0] _0896_;
  wire [2:0] _0897_;
  wire [2:0] _0898_;
  wire [2:0] _0899_;
  wire [2:0] _0900_;
  wire [2:0] _0901_;
  wire [2:0] _0902_;
  wire [2:0] _0903_;
  wire [2:0] _0904_;
  wire [2:0] _0905_;
  wire [2:0] _0906_;
  wire [2:0] _0907_;
  wire [2:0] _0908_;
  wire [2:0] _0909_;
  wire [2:0] _0910_;
  wire [2:0] _0911_;
  wire [2:0] _0912_;
  wire [2:0] _0913_;
  wire [2:0] _0914_;
  wire [2:0] _0915_;
  wire [2:0] _0916_;
  wire [2:0] _0917_;
  wire [2:0] _0918_;
  wire [31:0] _0919_;
  wire [31:0] _0920_;
  wire [31:0] _0921_;
  wire [31:0] _0922_;
  wire [31:0] _0923_;
  wire [31:0] _0924_;
  wire [31:0] _0925_;
  wire [31:0] _0926_;
  wire [31:0] _0927_;
  wire [31:0] _0928_;
  wire [31:0] _0929_;
  wire [31:0] _0930_;
  wire [31:0] _0931_;
  wire [31:0] _0932_;
  wire [31:0] _0933_;
  wire [31:0] _0934_;
  wire [31:0] _0935_;
  wire [31:0] _0936_;
  wire [31:0] _0937_;
  wire [31:0] _0938_;
  wire [31:0] _0939_;
  wire [31:0] _0940_;
  wire [31:0] _0941_;
  wire [31:0] _0942_;
  wire [31:0] _0943_;
  wire [31:0] _0944_;
  wire [31:0] _0945_;
  wire [31:0] _0946_;
  wire [31:0] _0947_;
  wire [31:0] _0948_;
  wire [31:0] _0949_;
  wire [31:0] _0950_;
  wire [31:0] _0951_;
  wire [31:0] _0952_;
  wire [31:0] _0953_;
  wire [31:0] _0954_;
  wire _0955_;
  wire _0956_;
  wire _0957_;
  wire _0958_;
  wire _0959_;
  wire _0960_;
  wire _0961_;
  wire _0962_;
  wire _0963_;
  wire _0964_;
  wire _0965_;
  wire _0966_;
  wire _0967_;
  wire _0968_;
  wire _0969_;
  wire _0970_;
  wire _0971_;
  wire _0972_;
  wire _0973_;
  wire _0974_;
  wire _0975_;
  wire _0976_;
  wire _0977_;
  wire _0978_;
  wire _0979_;
  wire _0980_;
  wire _0981_;
  wire _0982_;
  wire _0983_;
  wire _0984_;
  wire _0985_;
  wire _0986_;
  wire _0987_;
  wire _0988_;
  wire _0989_;
  wire _0990_;
  wire _0991_;
  wire _0992_;
  wire _0993_;
  wire _0994_;
  wire _0995_;
  wire _0996_;
  wire _0997_;
  wire _0998_;
  wire _0999_;
  wire _1000_;
  wire _1001_;
  wire _1002_;
  wire _1003_;
  wire _1004_;
  wire _1005_;
  wire _1006_;
  wire _1007_;
  wire _1008_;
  wire _1009_;
  wire _1010_;
  wire _1011_;
  wire _1012_;
  wire _1013_;
  wire _1014_;
  wire _1015_;
  wire _1016_;
  wire _1017_;
  wire _1018_;
  wire _1019_;
  wire _1020_;
  wire _1021_;
  wire _1022_;
  wire _1023_;
  wire _1024_;
  wire _1025_;
  wire _1026_;
  wire _1027_;
  wire _1028_;
  wire _1029_;
  wire _1030_;
  wire _1031_;
  wire _1032_;
  wire _1033_;
  wire _1034_;
  wire _1035_;
  wire _1036_;
  wire _1037_;
  wire _1038_;
  wire _1039_;
  wire _1040_;
  wire _1041_;
  wire _1042_;
  wire _1043_;
  wire _1044_;
  wire _1045_;
  wire _1046_;
  wire _1047_;
  wire _1048_;
  wire _1049_;
  wire _1050_;
  wire _1051_;
  wire _1052_;
  wire _1053_;
  wire _1054_;
  wire _1055_;
  wire _1056_;
  wire _1057_;
  wire _1058_;
  wire _1059_;
  wire _1060_;
  wire _1061_;
  wire _1062_;
  wire _1063_;
  wire _1064_;
  wire _1065_;
  wire _1066_;
  wire _1067_;
  wire _1068_;
  wire _1069_;
  wire _1070_;
  wire _1071_;
  wire _1072_;
  wire _1073_;
  wire _1074_;
  wire _1075_;
  wire _1076_;
  wire _1077_;
  wire _1078_;
  wire _1079_;
  wire _1080_;
  wire _1081_;
  wire _1082_;
  wire _1083_;
  wire _1084_;
  wire _1085_;
  wire _1086_;
  wire _1087_;
  wire _1088_;
  wire _1089_;
  wire _1090_;
  wire _1091_;
  wire _1092_;
  wire _1093_;
  wire _1094_;
  wire _1095_;
  wire _1096_;
  wire _1097_;
  wire _1098_;
  wire _1099_;
  wire _1100_;
  wire _1101_;
  wire _1102_;
  wire _1103_;
  wire _1104_;
  wire _1105_;
  wire _1106_;
  wire _1107_;
  wire _1108_;
  wire _1109_;
  wire _1110_;
  wire _1111_;
  wire [63:0] _1112_;
  wire [63:0] _1113_;
  wire [63:0] _1114_;
  wire [63:0] _1115_;
  wire [63:0] _1116_;
  wire [63:0] _1117_;
  wire [63:0] _1118_;
  wire [63:0] _1119_;
  wire [63:0] _1120_;
  wire [63:0] _1121_;
  wire [63:0] _1122_;
  wire [63:0] _1123_;
  wire [63:0] _1124_;
  wire [63:0] _1125_;
  wire [63:0] _1126_;
  wire [63:0] _1127_;
  wire [63:0] _1128_;
  wire [63:0] _1129_;
  wire [63:0] _1130_;
  wire [63:0] _1131_;
  wire [63:0] _1132_;
  wire [63:0] _1133_;
  wire [63:0] _1134_;
  wire [63:0] _1135_;
  wire [63:0] _1136_;
  wire [63:0] _1137_;
  wire [63:0] _1138_;
  wire [63:0] _1139_;
  wire [63:0] _1140_;
  wire [63:0] _1141_;
  wire [63:0] _1142_;
  wire [63:0] _1143_;
  wire [63:0] _1144_;
  wire [63:0] _1145_;
  wire [63:0] _1146_;
  wire [63:0] _1147_;
  wire [8:0] _1148_;
  wire [8:0] _1149_;
  wire [8:0] _1150_;
  wire [8:0] _1151_;
  wire [8:0] _1152_;
  wire [8:0] _1153_;
  wire [8:0] _1154_;
  wire [8:0] _1155_;
  wire [8:0] _1156_;
  wire [8:0] _1157_;
  wire [8:0] _1158_;
  wire [8:0] _1159_;
  wire [8:0] _1160_;
  wire [8:0] _1161_;
  wire [8:0] _1162_;
  wire [8:0] _1163_;
  wire [8:0] _1164_;
  wire [8:0] _1165_;
  wire [8:0] _1166_;
  wire [8:0] _1167_;
  wire [8:0] _1168_;
  wire [8:0] _1169_;
  wire [8:0] _1170_;
  wire [8:0] _1171_;
  wire [8:0] _1172_;
  wire [8:0] _1173_;
  wire [8:0] _1174_;
  wire [8:0] _1175_;
  wire [8:0] _1176_;
  wire [8:0] _1177_;
  wire [8:0] _1178_;
  wire [8:0] _1179_;
  wire [8:0] _1180_;
  wire [8:0] _1181_;
  wire [8:0] _1182_;
  wire [8:0] _1183_;
  wire [8:0] _1184_;
  wire [8:0] _1185_;
  wire [8:0] _1186_;
  wire [8:0] _1187_;
  wire [8:0] _1188_;
  wire [8:0] _1189_;
  wire [8:0] _1190_;
  wire [8:0] _1191_;
  wire [8:0] _1192_;
  wire [8:0] _1193_;
  wire [8:0] _1194_;
  wire [8:0] _1195_;
  wire [8:0] _1196_;
  wire [8:0] _1197_;
  wire [8:0] _1198_;
  wire [8:0] _1199_;
  wire [8:0] _1200_;
  wire [8:0] _1201_;
  wire [2:0] _1202_;
  wire [2:0] _1203_;
  wire [2:0] _1204_;
  wire [2:0] _1205_;
  wire [2:0] _1206_;
  wire [2:0] _1207_;
  wire [2:0] _1208_;
  wire [2:0] _1209_;
  wire [2:0] _1210_;
  wire [2:0] _1211_;
  wire [2:0] _1212_;
  wire [2:0] _1213_;
  wire [2:0] _1214_;
  wire [2:0] _1215_;
  wire [2:0] _1216_;
  wire [2:0] _1217_;
  wire [2:0] _1218_;
  wire [2:0] _1219_;
  wire [2:0] _1220_;
  wire [2:0] _1221_;
  wire [2:0] _1222_;
  wire [2:0] _1223_;
  wire [2:0] _1224_;
  wire [2:0] _1225_;
  wire [2:0] _1226_;
  wire [2:0] _1227_;
  wire [2:0] _1228_;
  wire [2:0] _1229_;
  wire [2:0] _1230_;
  wire [2:0] _1231_;
  wire [2:0] _1232_;
  wire [2:0] _1233_;
  wire [2:0] _1234_;
  wire [2:0] _1235_;
  wire [2:0] _1236_;
  wire [2:0] _1237_;
  wire [2:0] _1238_;
  wire [2:0] _1239_;
  wire [2:0] _1240_;
  wire [2:0] _1241_;
  wire [2:0] _1242_;
  wire [2:0] _1243_;
  wire [2:0] _1244_;
  wire [2:0] _1245_;
  wire [2:0] _1246_;
  wire [2:0] _1247_;
  wire [2:0] _1248_;
  wire [2:0] _1249_;
  wire [2:0] _1250_;
  wire [2:0] _1251_;
  wire [2:0] _1252_;
  wire [2:0] _1253_;
  wire [2:0] _1254_;
  wire [2:0] _1255_;
  wire [2:0] _1256_;
  wire [2:0] _1257_;
  wire [2:0] _1258_;
  wire [2:0] _1259_;
  wire [2:0] _1260_;
  wire [2:0] _1261_;
  wire [2:0] _1262_;
  wire [2:0] _1263_;
  wire [2:0] _1264_;
  wire [2:0] _1265_;
  wire [2:0] _1266_;
  wire [2:0] _1267_;
  wire [2:0] _1268_;
  wire [2:0] _1269_;
  wire [2:0] _1270_;
  wire [2:0] _1271_;
  wire [2:0] _1272_;
  wire [2:0] _1273_;
  wire [2:0] _1274_;
  wire [2:0] _1275_;
  wire [2:0] _1276_;
  wire [2:0] _1277_;
  wire [2:0] _1278_;
  wire [2:0] _1279_;
  wire [2:0] _1280_;
  wire [2:0] _1281_;
  wire [2:0] _1282_;
  wire [2:0] _1283_;
  wire [2:0] _1284_;
  wire [2:0] _1285_;
  wire [2:0] _1286_;
  wire [2:0] _1287_;
  wire [2:0] _1288_;
  wire [2:0] _1289_;
  wire [2:0] _1290_;
  wire [2:0] _1291_;
  wire [2:0] _1292_;
  wire _1293_;
  wire _1294_;
  wire _1295_;
  wire _1296_;
  wire _1297_;
  wire _1298_;
  wire _1299_;
  wire _1300_;
  wire _1301_;
  wire _1302_;
  wire _1303_;
  wire _1304_;
  wire _1305_;
  wire _1306_;
  wire _1307_;
  wire _1308_;
  wire _1309_;
  wire _1310_;
  wire _1311_;
  wire _1312_;
  wire _1313_;
  wire _1314_;
  wire _1315_;
  wire _1316_;
  wire _1317_;
  wire _1318_;
  wire _1319_;
  wire _1320_;
  wire _1321_;
  wire _1322_;
  wire _1323_;
  wire _1324_;
  wire _1325_;
  wire _1326_;
  wire _1327_;
  wire _1328_;
  wire _1329_;
  wire _1330_;
  wire _1331_;
  wire _1332_;
  wire _1333_;
  wire _1334_;
  wire _1335_;
  wire _1336_;
  wire _1337_;
  wire _1338_;
  wire _1339_;
  wire _1340_;
  wire _1341_;
  wire _1342_;
  wire _1343_;
  wire _1344_;
  wire _1345_;
  wire _1346_;
  wire _1347_;
  wire _1348_;
  wire _1349_;
  wire _1350_;
  wire _1351_;
  wire _1352_;
  wire _1353_;
  wire _1354_;
  wire _1355_;
  wire _1356_;
  wire _1357_;
  wire _1358_;
  wire _1359_;
  wire _1360_;
  wire _1361_;
  wire _1362_;
  wire _1363_;
  wire _1364_;
  wire _1365_;
  wire _1366_;
  wire _1367_;
  wire _1368_;
  wire _1369_;
  wire _1370_;
  wire _1371_;
  wire _1372_;
  wire _1373_;
  wire _1374_;
  wire _1375_;
  wire _1376_;
  wire _1377_;
  wire _1378_;
  wire _1379_;
  wire _1380_;
  wire _1381_;
  wire _1382_;
  wire _1383_;
  wire _1384_;
  wire _1385_;
  wire _1386_;
  wire _1387_;
  wire [2:0] _1388_;
  wire [2:0] _1389_;
  wire [2:0] _1390_;
  wire [2:0] _1391_;
  wire [2:0] _1392_;
  wire [2:0] _1393_;
  wire [2:0] _1394_;
  wire [2:0] _1395_;
  wire [2:0] _1396_;
  wire [2:0] _1397_;
  wire [2:0] _1398_;
  wire [2:0] _1399_;
  wire [2:0] _1400_;
  wire [2:0] _1401_;
  wire [2:0] _1402_;
  wire [2:0] _1403_;
  wire [2:0] _1404_;
  wire [2:0] _1405_;
  wire [2:0] _1406_;
  wire [2:0] _1407_;
  wire [2:0] _1408_;
  wire [2:0] _1409_;
  wire [2:0] _1410_;
  wire [2:0] _1411_;
  wire [2:0] _1412_;
  wire [2:0] _1413_;
  wire [2:0] _1414_;
  wire [2:0] _1415_;
  wire [2:0] _1416_;
  wire [2:0] _1417_;
  wire [2:0] _1418_;
  wire [2:0] _1419_;
  wire [2:0] _1420_;
  wire [2:0] _1421_;
  wire [2:0] _1422_;
  wire [2:0] _1423_;
  wire [2:0] _1424_;
  wire [2:0] _1425_;
  wire [2:0] _1426_;
  wire [2:0] _1427_;
  wire [2:0] _1428_;
  wire [2:0] _1429_;
  wire [2:0] _1430_;
  wire [2:0] _1431_;
  wire [2:0] _1432_;
  wire [2:0] _1433_;
  wire [2:0] _1434_;
  wire [2:0] _1435_;
  wire [2:0] _1436_;
  wire [2:0] _1437_;
  wire [2:0] _1438_;
  wire [2:0] _1439_;
  wire [2:0] _1440_;
  wire [2:0] _1441_;
  wire [2:0] _1442_;
  wire _1443_;
  wire _1444_;
  wire _1445_;
  wire _1446_;
  wire _1447_;
  wire _1448_;
  wire _1449_;
  wire _1450_;
  wire _1451_;
  wire _1452_;
  wire _1453_;
  wire _1454_;
  wire _1455_;
  wire _1456_;
  wire _1457_;
  wire _1458_;
  wire _1459_;
  wire _1460_;
  wire _1461_;
  wire _1462_;
  wire _1463_;
  wire _1464_;
  wire _1465_;
  wire _1466_;
  wire _1467_;
  wire _1468_;
  wire _1469_;
  wire _1470_;
  wire _1471_;
  wire _1472_;
  wire _1473_;
  wire _1474_;
  wire _1475_;
  wire _1476_;
  wire _1477_;
  wire _1478_;
  wire _1479_;
  wire _1480_;
  wire _1481_;
  wire _1482_;
  wire _1483_;
  wire _1484_;
  wire _1485_;
  wire _1486_;
  wire _1487_;
  wire _1488_;
  wire _1489_;
  wire _1490_;
  wire _1491_;
  wire _1492_;
  wire [1:0] _1493_;
  wire [1:0] _1494_;
  wire [31:0] _1495_;
  wire [31:0] _1496_;
  wire _1497_;
  wire _1498_;
  wire _1499_;
  wire _1500_;
  wire _1501_;
  wire _1502_;
  wire _1503_;
  wire _1504_;
  wire _1505_;
  wire _1506_;
  wire _1507_;
  wire _1508_;
  wire _1509_;
  wire _1510_;
  wire [30:0] _1511_;
  wire [1:0] _1512_;
  wire [1:0] _1513_;
  wire [1:0] _1514_;
  wire [1:0] _1515_;
  wire [31:0] _1516_;
  wire [31:0] _1517_;
  wire [31:0] _1518_;
  wire [31:0] _1519_;
  wire _1520_;
  wire _1521_;
  wire _1522_;
  wire _1523_;
  wire _1524_;
  wire _1525_;
  wire [31:0] _1526_;
  wire _1527_;
  wire _1528_;
  wire _1529_;
  wire _1530_;
  wire _1531_;
  wire _1532_;
  wire [1:0] _1533_;
  wire [1:0] _1534_;
  wire [1:0] _1535_;
  wire [1:0] _1536_;
  wire _1537_;
  wire _1538_;
  wire _1539_;
  wire _1540_;
  wire _1541_;
  wire _1542_;
  wire _1543_;
  wire _1544_;
  wire _1545_;
  wire _1546_;
  wire _1547_;
  wire [31:0] _1548_;
  wire [31:0] _1549_;
  wire [31:0] _1550_;
  wire _1551_;
  wire _1552_;
  wire [1:0] _1553_;
  wire [1:0] _1554_;
  wire [1:0] _1555_;
  wire _1556_;
  wire _1557_;
  wire [2:0] _1558_;
  wire [2:0] _1559_;
  wire [2:0] _1560_;
  wire [2:0] _1561_;
  wire [2:0] _1562_;
  wire [2:0] _1563_;
  wire [2:0] _1564_;
  wire [2:0] _1565_;
  wire [2:0] _1566_;
  wire [5:0] _1567_;
  wire [5:0] _1568_;
  wire [5:0] _1569_;
  wire [5:0] _1570_;
  wire [5:0] _1571_;
  wire [5:0] _1572_;
  wire _1573_;
  wire _1574_;
  wire [31:0] _1575_;
  wire [31:0] _1576_;
  wire [31:0] _1577_;
  wire _1578_;
  wire _1579_;
  wire [1:0] _1580_;
  wire [1:0] _1581_;
  wire [1:0] _1582_;
  wire _1583_;
  wire _1584_;
  wire _1585_;
  wire _1586_;
  wire _1587_;
  wire [31:0] _1588_;
  wire [31:0] _1589_;
  wire [31:0] _1590_;
  wire _1591_;
  wire _1592_;
  wire _1593_;
  wire _1594_;
  wire [31:0] _1595_;
  wire [31:0] _1596_;
  wire [31:0] _1597_;
  wire _1598_;
  wire _1599_;
  wire [2:0] _1600_;
  wire [2:0] _1601_;
  wire [2:0] _1602_;
  wire [1:0] _1603_;
  wire [1:0] _1604_;
  wire [1:0] _1605_;
  wire _1606_;
  wire _1607_;
  wire _1608_;
  wire _1609_;
  wire _1610_;
  wire [31:0] _1611_;
  wire [31:0] _1612_;
  wire [31:0] _1613_;
  wire _1614_;
  wire _1615_;
  wire _1616_;
  wire [5:0] _1617_;
  wire [5:0] _1618_;
  wire [5:0] _1619_;
  wire _1620_;
  wire _1621_;
  wire _1622_;
  wire [31:0] _1623_;
  wire [31:0] _1624_;
  wire [31:0] _1625_;
  wire _1626_;
  wire _1627_;
  wire _1628_;
  wire [3:0] _1629_;
  wire [3:0] _1630_;
  wire [3:0] _1631_;
  wire [31:0] _1632_;
  wire [31:0] _1633_;
  wire [31:0] _1634_;
  wire [31:0] _1635_;
  wire [31:0] _1636_;
  wire [31:0] _1637_;
  wire [31:0] _1638_;
  wire [31:0] _1639_;
  wire [31:0] _1640_;
  wire _1641_;
  wire _1642_;
  wire _1643_;
  wire _1644_;
  wire _1645_;
  wire [31:0] _1646_;
  wire [31:0] _1647_;
  wire [31:0] _1648_;
  wire _1649_;
  wire _1650_;
  wire _1651_;
  wire [2:0] _1652_;
  wire [2:0] _1653_;
  wire [2:0] _1654_;
  wire [1:0] _1655_;
  wire [1:0] _1656_;
  wire [1:0] _1657_;
  wire _1658_;
  wire _1659_;
  wire _1660_;
  wire [31:0] _1661_;
  wire [31:0] _1662_;
  wire [31:0] _1663_;
  wire _1664_;
  wire _1665_;
  wire _1666_;
  wire _1667_;
  wire _1668_;
  wire _1669_;
  wire _1670_;
  wire _1671_;
  wire _1672_;
  wire [5:0] _1673_;
  wire [5:0] _1674_;
  wire [5:0] _1675_;
  wire [5:0] _1676_;
  wire [5:0] _1677_;
  wire [5:0] _1678_;
  wire [5:0] _1679_;
  wire [5:0] _1680_;
  wire [5:0] _1681_;
  wire _1682_;
  wire _1683_;
  wire _1684_;
  wire _1685_;
  wire _1686_;
  wire _1687_;
  wire _1688_;
  wire _1689_;
  wire _1690_;
  wire [31:0] _1691_;
  wire [31:0] _1692_;
  wire [31:0] _1693_;
  wire [31:0] _1694_;
  wire [31:0] _1695_;
  wire [31:0] _1696_;
  wire [31:0] _1697_;
  wire [31:0] _1698_;
  wire [31:0] _1699_;
  wire _1700_;
  wire _1701_;
  wire _1702_;
  wire _1703_;
  wire _1704_;
  wire _1705_;
  wire _1706_;
  wire _1707_;
  wire _1708_;
  wire _1709_;
  wire [1:0] _1710_;
  wire [1:0] _1711_;
  wire [1:0] _1712_;
  wire [1:0] _1713_;
  wire [1:0] _1714_;
  wire [1:0] _1715_;
  wire [1:0] _1716_;
  wire [1:0] _1717_;
  wire [1:0] _1718_;
  wire [3:0] _1719_;
  wire [3:0] _1720_;
  wire [3:0] _1721_;
  wire [1:0] _1722_;
  wire [1:0] _1723_;
  wire [1:0] _1724_;
  wire [1:0] _1725_;
  wire [1:0] _1726_;
  wire [1:0] _1727_;
  wire _1728_;
  wire _1729_;
  wire _1730_;
  wire _1731_;
  wire _1732_;
  wire [11:0] _1733_;
  wire [11:0] _1734_;
  wire [11:0] _1735_;
  wire [1:0] _1736_;
  wire [1:0] _1737_;
  wire [1:0] _1738_;
  wire [1:0] _1739_;
  wire [1:0] _1740_;
  wire [1:0] _1741_;
  wire _1742_;
  wire _1743_;
  wire _1744_;
  wire _1745_;
  wire _1746_;
  wire _1747_;
  wire _1748_;
  wire _1749_;
  wire _1750_;
  wire [1:0] _1751_;
  wire [1:0] _1752_;
  wire [1:0] _1753_;
  wire _1754_;
  wire _1755_;
  wire [1:0] _1756_;
  wire [1:0] _1757_;
  wire [1:0] _1758_;
  wire _1759_;
  wire _1760_;
  wire [1:0] _1761_;
  wire [1:0] _1762_;
  wire [1:0] _1763_;
  wire [31:0] _1764_;
  wire [31:0] _1765_;
  wire [31:0] _1766_;
  wire [31:0] _1767_;
  wire [31:0] _1768_;
  wire [31:0] _1769_;
  wire _1770_;
  wire _1771_;
  wire _1772_;
  wire _1773_;
  wire _1774_;
  wire _1775_;
  wire [31:0] _1776_;
  wire [31:0] _1777_;
  wire [31:0] _1778_;
  wire [31:0] _1779_;
  wire [31:0] _1780_;
  wire _1781_;
  wire _1782_;
  wire _1783_;
  wire _1784_;
  wire _1785_;
  wire _1786_;
  wire _1787_;
  wire _1788_;
  wire _1789_;
  wire _1790_;
  wire [31:0] _1791_;
  wire [31:0] _1792_;
  wire [31:0] _1793_;
  wire _1794_;
  wire _1795_;
  wire _1796_;
  wire _1797_;
  wire _1798_;
  wire _1799_;
  wire _1800_;
  wire _1801_;
  wire _1802_;
  wire _1803_;
  wire _1804_;
  wire _1805_;
  wire _1806_;
  wire _1807_;
  wire _1808_;
  wire [5:0] _1809_;
  wire [5:0] _1810_;
  wire [5:0] _1811_;
  wire [30:0] _1812_;
  wire [28:0] _1813_;
  wire [11:0] _1814_;
  wire [11:0] _1815_;
  wire [11:0] _1816_;
  wire [4:0] _1817_;
  wire [4:0] _1818_;
  wire [4:0] _1819_;
  wire [4:0] _1820_;
  wire [4:0] _1821_;
  wire [4:0] _1822_;
  wire [4:0] _1823_;
  wire [4:0] _1824_;
  wire [4:0] _1825_;
  wire [4:0] _1826_;
  wire [4:0] _1827_;
  wire [4:0] _1828_;
  wire [4:0] _1829_;
  wire [4:0] _1830_;
  wire [4:0] _1831_;
  wire [4:0] _1832_;
  wire [4:0] _1833_;
  wire [4:0] _1834_;
  wire [4:0] _1835_;
  wire [4:0] _1836_;
  wire [4:0] _1837_;
  wire [4:0] _1838_;
  wire [4:0] _1839_;
  wire [4:0] _1840_;
  wire [4:0] _1841_;
  wire [4:0] _1842_;
  wire [4:0] _1843_;
  wire [4:0] _1844_;
  wire [4:0] _1845_;
  wire [4:0] _1846_;
  wire [4:0] _1847_;
  wire [4:0] _1848_;
  wire [11:0] _1849_;
  wire [11:0] _1850_;
  wire [11:0] _1851_;
  wire [11:0] _1852_;
  wire [11:0] _1853_;
  wire [11:0] _1854_;
  wire [11:0] _1855_;
  wire [11:0] _1856_;
  wire [11:0] _1857_;
  wire [11:0] _1858_;
  wire [11:0] _1859_;
  wire [11:0] _1860_;
  wire [11:0] _1861_;
  wire [11:0] _1862_;
  wire [11:0] _1863_;
  wire [11:0] _1864_;
  wire [11:0] _1865_;
  wire [11:0] _1866_;
  wire [11:0] _1867_;
  wire [11:0] _1868_;
  wire [11:0] _1869_;
  wire [11:0] _1870_;
  wire [11:0] _1871_;
  wire [11:0] _1872_;
  wire [11:0] _1873_;
  wire [11:0] _1874_;
  wire [11:0] _1875_;
  wire [11:0] _1876_;
  wire [11:0] _1877_;
  wire [11:0] _1878_;
  wire [11:0] _1879_;
  wire [11:0] _1880_;
  wire [11:0] _1881_;
  wire [30:0] _1882_;
  wire [11:0] _1883_;
  wire [11:0] _1884_;
  wire [11:0] _1885_;
  wire [11:0] _1886_;
  wire [11:0] _1887_;
  wire [11:0] _1888_;
  wire [11:0] _1889_;
  wire [11:0] _1890_;
  wire [11:0] _1891_;
  wire [11:0] _1892_;
  wire [11:0] _1893_;
  wire [11:0] _1894_;
  wire [11:0] _1895_;
  wire [11:0] _1896_;
  wire [11:0] _1897_;
  wire [11:0] _1898_;
  wire [11:0] _1899_;
  wire [11:0] _1900_;
  wire [11:0] _1901_;
  wire [11:0] _1902_;
  wire [11:0] _1903_;
  wire [11:0] _1904_;
  wire [11:0] _1905_;
  wire [11:0] _1906_;
  wire [11:0] _1907_;
  wire [11:0] _1908_;
  wire [11:0] _1909_;
  wire [11:0] _1910_;
  wire [11:0] _1911_;
  wire [11:0] _1912_;
  wire [11:0] _1913_;
  wire [11:0] _1914_;
  wire [11:0] _1915_;
  wire [11:0] _1916_;
  wire [11:0] _1917_;
  wire [11:0] _1918_;
  wire [11:0] _1919_;
  wire [11:0] _1920_;
  wire [11:0] _1921_;
  wire [11:0] _1922_;
  wire [11:0] _1923_;
  wire [11:0] _1924_;
  wire [11:0] _1925_;
  wire [11:0] _1926_;
  wire [11:0] _1927_;
  wire [11:0] _1928_;
  wire [11:0] _1929_;
  wire [11:0] _1930_;
  wire [11:0] _1931_;
  wire [11:0] _1932_;
  wire [11:0] _1933_;
  wire [11:0] _1934_;
  wire [11:0] _1935_;
  wire [11:0] _1936_;
  wire [11:0] _1937_;
  wire [11:0] _1938_;
  wire [11:0] _1939_;
  wire [11:0] _1940_;
  wire [11:0] _1941_;
  wire [11:0] _1942_;
  wire [11:0] _1943_;
  wire [11:0] _1944_;
  wire [11:0] _1945_;
  wire [11:0] _1946_;
  wire [11:0] _1947_;
  wire [11:0] _1948_;
  wire [11:0] _1949_;
  wire [11:0] _1950_;
  wire [11:0] _1951_;
  wire [11:0] _1952_;
  wire [11:0] _1953_;
  wire [11:0] _1954_;
  wire [11:0] _1955_;
  wire [11:0] _1956_;
  wire [11:0] _1957_;
  wire [11:0] _1958_;
  wire [11:0] _1959_;
  wire [11:0] _1960_;
  wire [11:0] _1961_;
  wire [11:0] _1962_;
  wire [11:0] _1963_;
  wire [11:0] _1964_;
  wire [11:0] _1965_;
  wire [11:0] _1966_;
  wire [11:0] _1967_;
  wire [11:0] _1968_;
  wire [11:0] _1969_;
  wire [11:0] _1970_;
  wire [11:0] _1971_;
  wire [11:0] _1972_;
  wire [11:0] _1973_;
  wire [11:0] _1974_;
  wire [11:0] _1975_;
  wire [11:0] _1976_;
  wire [11:0] _1977_;
  wire [11:0] _1978_;
  wire [11:0] _1979_;
  wire [11:0] _1980_;
  wire [11:0] _1981_;
  wire [11:0] _1982_;
  wire [2:0] _1983_;
  wire [17:0] _1984_;
  wire [31:0] _1985_;
  wire [31:0] _1986_;
  wire [31:0] _1987_;
  wire [1:0] _1988_;
  wire [1:0] _1989_;
  wire [1:0] _1990_;
  wire _1991_;
  wire _1992_;
  wire _1993_;
  wire _1994_;
  wire _1995_;
  wire _1996_;
  wire _1997_;
  wire _1998_;
  wire _1999_;
  wire _2000_;
  wire _2001_;
  wire _2002_;
  wire _2003_;
  wire _2004_;
  wire _2005_;
  wire _2006_;
  wire _2007_;
  wire _2008_;
  wire _2009_;
  wire _2010_;
  wire _2011_;
  wire _2012_;
  wire _2013_;
  wire _2014_;
  wire _2015_;
  wire _2016_;
  wire _2017_;
  wire _2018_;
  wire _2019_;
  wire _2020_;
  wire _2021_;
  wire _2022_;
  wire _2023_;
  wire _2024_;
  wire [31:0] _2025_;
  wire _2026_;
  wire [31:0] _2027_;
  wire _2028_;
  wire _2029_;
  wire [17:0] _2030_;
  wire _2031_;
  wire _2032_;
  wire _2033_;
  wire _2034_;
  wire _2035_;
  wire _2036_;
  wire _2037_;
  wire _2038_;
  wire _2039_;
  wire _2040_;
  wire _2041_;
  wire _2042_;
  wire _2043_;
  wire _2044_;
  wire _2045_;
  wire _2046_;
  wire _2047_;
  wire _2048_;
  wire [11:0] _2049_;
  wire [11:0] _2050_;
  wire [11:0] _2051_;
  wire [11:0] _2052_;
  wire _2053_;
  wire _2054_;
  wire _2055_;
  wire _2056_;
  wire _2057_;
  wire _2058_;
  wire _2059_;
  wire _2060_;
  wire _2061_;
  wire _2062_;
  wire _2063_;
  wire _2064_;
  wire _2065_;
  wire _2066_;
  wire _2067_;
  wire _2068_;
  wire [31:0] _2069_;
  wire [31:0] _2070_;
  wire [31:0] _2071_;
  wire [31:0] _2072_;
  wire [31:0] _2073_;
  wire [31:0] _2074_;
  wire _2075_;
  wire _2076_;
  wire _2077_;
  wire _2078_;
  wire _2079_;
  wire _2080_;
  wire _2081_;
  wire _2082_;
  wire _2083_;
  wire _2084_;
  wire _2085_;
  wire _2086_;
  wire _2087_;
  wire _2088_;
  wire _2089_;
  wire _2090_;
  wire _2091_;
  wire _2092_;
  wire _2093_;
  wire _2094_;
  wire _2095_;
  wire _2096_;
  wire _2097_;
  wire _2098_;
  wire _2099_;
  wire _2100_;
  wire _2101_;
  wire _2102_;
  wire _2103_;
  wire _2104_;
  wire _2105_;
  wire _2106_;
  wire _2107_;
  wire _2108_;
  wire _2109_;
  wire _2110_;
  wire _2111_;
  wire _2112_;
  wire _2113_;
  wire _2114_;
  wire _2115_;
  wire _2116_;
  wire [2:0] _2117_;
  wire [2:0] _2118_;
  wire [2:0] _2119_;
  wire [2:0] _2120_;
  wire [2:0] _2121_;
  wire [2:0] _2122_;
  wire [2:0] _2123_;
  wire [2:0] _2124_;
  wire [2:0] _2125_;
  wire [2:0] _2126_;
  wire [2:0] _2127_;
  wire [2:0] _2128_;
  wire [2:0] _2129_;
  wire [2:0] _2130_;
  wire [2:0] _2131_;
  wire [2:0] _2132_;
  wire [2:0] _2133_;
  wire [2:0] _2134_;
  wire [2:0] _2135_;
  wire [2:0] _2136_;
  wire [2:0] _2137_;
  wire [2:0] _2138_;
  wire [2:0] _2139_;
  wire [2:0] _2140_;
  wire [2:0] _2141_;
  wire [2:0] _2142_;
  wire [2:0] _2143_;
  wire [2:0] _2144_;
  wire [2:0] _2145_;
  wire [2:0] _2146_;
  wire [2:0] _2147_;
  wire [2:0] _2148_;
  wire [2:0] _2149_;
  wire [2:0] _2150_;
  wire [2:0] _2151_;
  wire [2:0] _2152_;
  wire [2:0] _2153_;
  wire [2:0] _2154_;
  wire [2:0] _2155_;
  wire [2:0] _2156_;
  wire [2:0] _2157_;
  wire [2:0] _2158_;
  wire [2:0] _2159_;
  wire [2:0] _2160_;
  wire [2:0] _2161_;
  wire _2162_;
  wire _2163_;
  wire _2164_;
  wire _2165_;
  wire _2166_;
  wire _2167_;
  wire _2168_;
  wire _2169_;
  wire _2170_;
  wire _2171_;
  wire _2172_;
  wire _2173_;
  wire _2174_;
  wire _2175_;
  wire _2176_;
  wire _2177_;
  wire _2178_;
  wire _2179_;
  wire _2180_;
  wire _2181_;
  wire _2182_;
  wire _2183_;
  wire _2184_;
  wire _2185_;
  wire _2186_;
  wire _2187_;
  wire _2188_;
  wire _2189_;
  wire _2190_;
  wire _2191_;
  wire _2192_;
  wire _2193_;
  wire _2194_;
  wire _2195_;
  wire [2:0] _2196_;
  wire [2:0] _2197_;
  wire [2:0] _2198_;
  wire [2:0] _2199_;
  wire [2:0] _2200_;
  wire [2:0] _2201_;
  wire [2:0] _2202_;
  wire [2:0] _2203_;
  wire [2:0] _2204_;
  wire [2:0] _2205_;
  wire [2:0] _2206_;
  wire [2:0] _2207_;
  wire [2:0] _2208_;
  wire [2:0] _2209_;
  wire [2:0] _2210_;
  wire [2:0] _2211_;
  wire [2:0] _2212_;
  wire [2:0] _2213_;
  wire [2:0] _2214_;
  wire [2:0] _2215_;
  wire [2:0] _2216_;
  wire [2:0] _2217_;
  wire [2:0] _2218_;
  wire [2:0] _2219_;
  wire [2:0] _2220_;
  wire [2:0] _2221_;
  wire [2:0] _2222_;
  wire [2:0] _2223_;
  wire [2:0] _2224_;
  wire [2:0] _2225_;
  wire [2:0] _2226_;
  wire [2:0] _2227_;
  wire [2:0] _2228_;
  wire [2:0] _2229_;
  wire [2:0] _2230_;
  wire [2:0] _2231_;
  wire [2:0] _2232_;
  wire [2:0] _2233_;
  wire [2:0] _2234_;
  wire [2:0] _2235_;
  wire [2:0] _2236_;
  wire [31:0] _2237_;
  wire [31:0] _2238_;
  wire [31:0] _2239_;
  wire [31:0] _2240_;
  wire [31:0] _2241_;
  wire [31:0] _2242_;
  wire [31:0] _2243_;
  wire [31:0] _2244_;
  wire [31:0] _2245_;
  wire [31:0] _2246_;
  wire [31:0] _2247_;
  wire [31:0] _2248_;
  wire [31:0] _2249_;
  wire [31:0] _2250_;
  wire [31:0] _2251_;
  wire [31:0] _2252_;
  wire [31:0] _2253_;
  wire [31:0] _2254_;
  wire [31:0] _2255_;
  wire [31:0] _2256_;
  wire [31:0] _2257_;
  wire [31:0] _2258_;
  wire [31:0] _2259_;
  wire [31:0] _2260_;
  wire [31:0] _2261_;
  wire [31:0] _2262_;
  wire [31:0] _2263_;
  wire [31:0] _2264_;
  wire [31:0] _2265_;
  wire [31:0] _2266_;
  wire [31:0] _2267_;
  wire [31:0] _2268_;
  wire [31:0] _2269_;
  wire [31:0] _2270_;
  wire [31:0] _2271_;
  wire [31:0] _2272_;
  wire _2273_;
  wire _2274_;
  wire _2275_;
  wire _2276_;
  wire _2277_;
  wire _2278_;
  wire _2279_;
  wire _2280_;
  wire _2281_;
  wire _2282_;
  wire _2283_;
  wire _2284_;
  wire _2285_;
  wire _2286_;
  wire _2287_;
  wire _2288_;
  wire _2289_;
  wire _2290_;
  wire _2291_;
  wire _2292_;
  wire _2293_;
  wire _2294_;
  wire _2295_;
  wire _2296_;
  wire _2297_;
  wire _2298_;
  wire _2299_;
  wire _2300_;
  wire _2301_;
  wire _2302_;
  wire _2303_;
  wire _2304_;
  wire _2305_;
  wire _2306_;
  wire _2307_;
  wire _2308_;
  wire _2309_;
  wire _2310_;
  wire _2311_;
  wire _2312_;
  wire _2313_;
  wire _2314_;
  wire _2315_;
  wire _2316_;
  wire _2317_;
  wire _2318_;
  wire _2319_;
  wire _2320_;
  wire _2321_;
  wire _2322_;
  wire _2323_;
  wire _2324_;
  wire _2325_;
  wire _2326_;
  wire _2327_;
  wire _2328_;
  wire _2329_;
  wire _2330_;
  wire _2331_;
  wire _2332_;
  wire _2333_;
  wire _2334_;
  wire _2335_;
  wire _2336_;
  wire _2337_;
  wire _2338_;
  wire _2339_;
  wire _2340_;
  wire _2341_;
  wire _2342_;
  wire _2343_;
  wire _2344_;
  wire _2345_;
  wire _2346_;
  wire [63:0] _2347_;
  wire [63:0] _2348_;
  wire [63:0] _2349_;
  wire [63:0] _2350_;
  wire [63:0] _2351_;
  wire [63:0] _2352_;
  wire [63:0] _2353_;
  wire [63:0] _2354_;
  wire [63:0] _2355_;
  wire [63:0] _2356_;
  wire [63:0] _2357_;
  wire [63:0] _2358_;
  wire [63:0] _2359_;
  wire [63:0] _2360_;
  wire [63:0] _2361_;
  wire [63:0] _2362_;
  wire [63:0] _2363_;
  wire [63:0] _2364_;
  wire [63:0] _2365_;
  wire [63:0] _2366_;
  wire [63:0] _2367_;
  wire [63:0] _2368_;
  wire [63:0] _2369_;
  wire [63:0] _2370_;
  wire [63:0] _2371_;
  wire [63:0] _2372_;
  wire [63:0] _2373_;
  wire [63:0] _2374_;
  wire [63:0] _2375_;
  wire [63:0] _2376_;
  wire [63:0] _2377_;
  wire [63:0] _2378_;
  wire [63:0] _2379_;
  wire [63:0] _2380_;
  wire [63:0] _2381_;
  wire [63:0] _2382_;
  wire [8:0] _2383_;
  wire [8:0] _2384_;
  wire [8:0] _2385_;
  wire [8:0] _2386_;
  wire [8:0] _2387_;
  wire [8:0] _2388_;
  wire [8:0] _2389_;
  wire [8:0] _2390_;
  wire [8:0] _2391_;
  wire [8:0] _2392_;
  wire [8:0] _2393_;
  wire [8:0] _2394_;
  wire [8:0] _2395_;
  wire [8:0] _2396_;
  wire [8:0] _2397_;
  wire [8:0] _2398_;
  wire [8:0] _2399_;
  wire [8:0] _2400_;
  wire [8:0] _2401_;
  wire [8:0] _2402_;
  wire [8:0] _2403_;
  wire [8:0] _2404_;
  wire [8:0] _2405_;
  wire [8:0] _2406_;
  wire [8:0] _2407_;
  wire [8:0] _2408_;
  wire [8:0] _2409_;
  wire [8:0] _2410_;
  wire [8:0] _2411_;
  wire [8:0] _2412_;
  wire [8:0] _2413_;
  wire [8:0] _2414_;
  wire [8:0] _2415_;
  wire [8:0] _2416_;
  wire [8:0] _2417_;
  wire [8:0] _2418_;
  wire [8:0] _2419_;
  wire [8:0] _2420_;
  wire [8:0] _2421_;
  wire [8:0] _2422_;
  wire [8:0] _2423_;
  wire [8:0] _2424_;
  wire [8:0] _2425_;
  wire [8:0] _2426_;
  wire [8:0] _2427_;
  wire [8:0] _2428_;
  wire [8:0] _2429_;
  wire [8:0] _2430_;
  wire [8:0] _2431_;
  wire [8:0] _2432_;
  wire [8:0] _2433_;
  wire [8:0] _2434_;
  wire [8:0] _2435_;
  wire [8:0] _2436_;
  wire [2:0] _2437_;
  wire [2:0] _2438_;
  wire [2:0] _2439_;
  wire [2:0] _2440_;
  wire [2:0] _2441_;
  wire [2:0] _2442_;
  wire [2:0] _2443_;
  wire [2:0] _2444_;
  wire [2:0] _2445_;
  wire [2:0] _2446_;
  wire [2:0] _2447_;
  wire [2:0] _2448_;
  wire [2:0] _2449_;
  wire [2:0] _2450_;
  wire [2:0] _2451_;
  wire [2:0] _2452_;
  wire [2:0] _2453_;
  wire [2:0] _2454_;
  wire [2:0] _2455_;
  wire [2:0] _2456_;
  wire [2:0] _2457_;
  wire [2:0] _2458_;
  wire [2:0] _2459_;
  wire [2:0] _2460_;
  wire [2:0] _2461_;
  wire [2:0] _2462_;
  wire [2:0] _2463_;
  wire [2:0] _2464_;
  wire [2:0] _2465_;
  wire [2:0] _2466_;
  wire [2:0] _2467_;
  wire [2:0] _2468_;
  wire [2:0] _2469_;
  wire [2:0] _2470_;
  wire [2:0] _2471_;
  wire [2:0] _2472_;
  wire [2:0] _2473_;
  wire [2:0] _2474_;
  wire [2:0] _2475_;
  wire [2:0] _2476_;
  wire [2:0] _2477_;
  wire [2:0] _2478_;
  wire [2:0] _2479_;
  wire [2:0] _2480_;
  wire [2:0] _2481_;
  wire [2:0] _2482_;
  wire [2:0] _2483_;
  wire [2:0] _2484_;
  wire [2:0] _2485_;
  wire [2:0] _2486_;
  wire [2:0] _2487_;
  wire [2:0] _2488_;
  wire [2:0] _2489_;
  wire [2:0] _2490_;
  wire [2:0] _2491_;
  wire [2:0] _2492_;
  wire [2:0] _2493_;
  wire [2:0] _2494_;
  wire [2:0] _2495_;
  wire _2496_;
  wire _2497_;
  wire _2498_;
  wire _2499_;
  wire _2500_;
  wire _2501_;
  wire _2502_;
  wire _2503_;
  wire _2504_;
  wire _2505_;
  wire _2506_;
  wire _2507_;
  wire _2508_;
  wire _2509_;
  wire _2510_;
  wire _2511_;
  wire _2512_;
  wire _2513_;
  wire _2514_;
  wire _2515_;
  wire _2516_;
  wire _2517_;
  wire _2518_;
  wire _2519_;
  wire _2520_;
  wire _2521_;
  wire _2522_;
  wire _2523_;
  wire _2524_;
  wire _2525_;
  wire _2526_;
  wire _2527_;
  wire _2528_;
  wire [2:0] _2529_;
  wire [2:0] _2530_;
  wire [2:0] _2531_;
  wire [2:0] _2532_;
  wire [2:0] _2533_;
  wire [2:0] _2534_;
  wire [2:0] _2535_;
  wire [2:0] _2536_;
  wire [2:0] _2537_;
  wire [2:0] _2538_;
  wire [2:0] _2539_;
  wire [2:0] _2540_;
  wire [2:0] _2541_;
  wire [2:0] _2542_;
  wire [2:0] _2543_;
  wire [2:0] _2544_;
  wire [2:0] _2545_;
  wire [2:0] _2546_;
  wire [2:0] _2547_;
  wire [2:0] _2548_;
  wire [2:0] _2549_;
  wire [2:0] _2550_;
  wire [2:0] _2551_;
  wire [2:0] _2552_;
  wire [2:0] _2553_;
  wire [2:0] _2554_;
  wire [2:0] _2555_;
  wire [2:0] _2556_;
  wire [2:0] _2557_;
  wire _2558_;
  wire _2559_;
  wire _2560_;
  wire _2561_;
  wire _2562_;
  wire _2563_;
  wire _2564_;
  wire _2565_;
  wire _2566_;
  wire _2567_;
  wire _2568_;
  wire _2569_;
  wire _2570_;
  wire _2571_;
  wire _2572_;
  wire _2573_;
  wire _2574_;
  wire _2575_;
  wire _2576_;
  wire _2577_;
  wire _2578_;
  wire _2579_;
  wire _2580_;
  wire _2581_;
  wire _2582_;
  wire _2583_;
  wire [31:0] _2584_;
  wire _2585_;
  wire _2586_;
  wire _2587_;
  wire _2588_;
  wire _2589_;
  wire _2590_;
  wire _2591_;
  wire _2592_;
  wire [30:0] _2593_;
  wire [31:0] _2594_;
  wire [31:0] _2595_;
  wire _2596_;
  wire _2597_;
  wire [31:0] _2598_;
  wire _2599_;
  wire _2600_;
  wire _2601_;
  wire _2602_;
  wire _2603_;
  wire _2604_;
  wire _2605_;
  wire _2606_;
  wire _2607_;
  wire _2608_;
  wire _2609_;
  wire _2610_;
  wire _2611_;
  wire [31:0] _2612_;
  wire [31:0] _2613_;
  wire [31:0] _2614_;
  wire [1:0] _2615_;
  wire [1:0] _2616_;
  wire [1:0] _2617_;
  wire [2:0] _2618_;
  wire [2:0] _2619_;
  wire [2:0] _2620_;
  wire [2:0] _2621_;
  wire [2:0] _2622_;
  wire [2:0] _2623_;
  wire [2:0] _2624_;
  wire [2:0] _2625_;
  wire [2:0] _2626_;
  wire [5:0] _2627_;
  wire [5:0] _2628_;
  wire [5:0] _2629_;
  wire [5:0] _2630_;
  wire [5:0] _2631_;
  wire [5:0] _2632_;
  wire _2633_;
  wire _2634_;
  wire [31:0] _2635_;
  wire [31:0] _2636_;
  wire [31:0] _2637_;
  wire [1:0] _2638_;
  wire [1:0] _2639_;
  wire [1:0] _2640_;
  wire _2641_;
  wire [31:0] _2642_;
  wire _2643_;
  wire _2644_;
  wire [31:0] _2645_;
  wire [31:0] _2646_;
  wire [31:0] _2647_;
  wire [2:0] _2648_;
  wire [2:0] _2649_;
  wire [2:0] _2650_;
  wire [1:0] _2651_;
  wire [1:0] _2652_;
  wire [1:0] _2653_;
  wire _2654_;
  wire [31:0] _2655_;
  wire _2656_;
  wire [5:0] _2657_;
  wire [5:0] _2658_;
  wire [5:0] _2659_;
  wire _2660_;
  wire [31:0] _2661_;
  wire _2662_;
  wire [3:0] _2663_;
  wire [3:0] _2664_;
  wire [3:0] _2665_;
  wire [31:0] _2666_;
  wire [31:0] _2667_;
  wire [31:0] _2668_;
  wire [31:0] _2669_;
  wire [31:0] _2670_;
  wire [31:0] _2671_;
  wire [31:0] _2672_;
  wire [31:0] _2673_;
  wire [31:0] _2674_;
  wire _2675_;
  wire [31:0] _2676_;
  wire [31:0] _2677_;
  wire [31:0] _2678_;
  wire _2679_;
  wire [2:0] _2680_;
  wire [1:0] _2681_;
  wire [1:0] _2682_;
  wire [1:0] _2683_;
  wire _2684_;
  wire [31:0] _2685_;
  wire _2686_;
  wire _2687_;
  wire _2688_;
  wire [5:0] _2689_;
  wire [5:0] _2690_;
  wire [5:0] _2691_;
  wire [5:0] _2692_;
  wire [5:0] _2693_;
  wire [5:0] _2694_;
  wire [5:0] _2695_;
  wire [5:0] _2696_;
  wire [5:0] _2697_;
  wire _2698_;
  wire _2699_;
  wire _2700_;
  wire [31:0] _2701_;
  wire [31:0] _2702_;
  wire [31:0] _2703_;
  wire [31:0] _2704_;
  wire [31:0] _2705_;
  wire [31:0] _2706_;
  wire [31:0] _2707_;
  wire _2708_;
  wire _2709_;
  wire [1:0] _2710_;
  wire [1:0] _2711_;
  wire [1:0] _2712_;
  wire [1:0] _2713_;
  wire [1:0] _2714_;
  wire [1:0] _2715_;
  wire [1:0] _2716_;
  wire [3:0] _2717_;
  wire [3:0] _2718_;
  wire [3:0] _2719_;
  wire [1:0] _2720_;
  wire [1:0] _2721_;
  wire [1:0] _2722_;
  wire [1:0] _2723_;
  wire _2724_;
  wire [11:0] _2725_;
  wire [11:0] _2726_;
  wire [11:0] _2727_;
  wire [1:0] _2728_;
  wire [1:0] _2729_;
  wire [1:0] _2730_;
  wire [1:0] _2731_;
  wire _2732_;
  wire [1:0] _2733_;
  wire [1:0] _2734_;
  wire [1:0] _2735_;
  wire [1:0] _2736_;
  wire [1:0] _2737_;
  wire [1:0] _2738_;
  wire [1:0] _2739_;
  wire [31:0] _2740_;
  wire [31:0] _2741_;
  wire [31:0] _2742_;
  wire [31:0] _2743_;
  wire [31:0] _2744_;
  wire [31:0] _2745_;
  wire _2746_;
  wire _2747_;
  wire [31:0] _2748_;
  wire [31:0] _2749_;
  wire [31:0] _2750_;
  wire [31:0] _2751_;
  wire [31:0] _2752_;
  wire _2753_;
  wire [5:0] _2754_;
  wire [5:0] _2755_;
  wire [5:0] _2756_;
  wire [31:0] _2757_;
  wire [31:0] _2758_;
  wire [31:0] _2759_;
  wire [1:0] _2760_;
  wire [1:0] _2761_;
  wire [1:0] _2762_;
  wire _2763_;
  wire [11:0] _2764_;
  wire [31:0] _2765_;
  wire [31:0] _2766_;
  wire _2767_;
  wire _2768_;
  wire _2769_;
  wire _2770_;
  wire _2771_;
  wire _2772_;
  wire _2773_;
  wire _2774_;
  wire _2775_;
  wire _2776_;
  wire _2777_;
  wire _2778_;
  wire _2779_;
  wire [2:0] _2780_;
  wire [2:0] _2781_;
  wire [2:0] _2782_;
  wire [2:0] _2783_;
  wire [2:0] _2784_;
  wire [2:0] _2785_;
  wire [2:0] _2786_;
  wire [2:0] _2787_;
  wire [2:0] _2788_;
  wire [2:0] _2789_;
  wire [2:0] _2790_;
  wire [2:0] _2791_;
  wire [2:0] _2792_;
  wire [2:0] _2793_;
  wire _2794_;
  wire _2795_;
  wire _2796_;
  wire _2797_;
  wire _2798_;
  wire _2799_;
  wire _2800_;
  wire _2801_;
  wire _2802_;
  wire _2803_;
  wire _2804_;
  wire _2805_;
  wire _2806_;
  wire _2807_;
  wire _2808_;
  wire _2809_;
  wire [2:0] _2810_;
  wire [2:0] _2811_;
  wire [2:0] _2812_;
  wire [2:0] _2813_;
  wire [2:0] _2814_;
  wire [2:0] _2815_;
  wire [2:0] _2816_;
  wire [2:0] _2817_;
  wire [2:0] _2818_;
  wire [2:0] _2819_;
  wire [2:0] _2820_;
  wire [2:0] _2821_;
  wire [2:0] _2822_;
  wire [2:0] _2823_;
  wire [2:0] _2824_;
  wire [2:0] _2825_;
  wire [31:0] _2826_;
  wire [31:0] _2827_;
  wire [31:0] _2828_;
  wire [31:0] _2829_;
  wire [31:0] _2830_;
  wire [31:0] _2831_;
  wire [31:0] _2832_;
  wire _2833_;
  wire _2834_;
  wire _2835_;
  wire _2836_;
  wire _2837_;
  wire _2838_;
  wire _2839_;
  wire _2840_;
  wire _2841_;
  wire _2842_;
  wire _2843_;
  wire _2844_;
  wire _2845_;
  wire _2846_;
  wire _2847_;
  wire _2848_;
  wire _2849_;
  wire _2850_;
  wire _2851_;
  wire _2852_;
  wire _2853_;
  wire _2854_;
  wire _2855_;
  wire _2856_;
  wire _2857_;
  wire _2858_;
  wire _2859_;
  wire _2860_;
  wire _2861_;
  wire _2862_;
  wire _2863_;
  wire _2864_;
  wire _2865_;
  wire _2866_;
  wire _2867_;
  wire _2868_;
  wire _2869_;
  wire _2870_;
  wire _2871_;
  wire _2872_;
  wire _2873_;
  wire _2874_;
  wire _2875_;
  wire _2876_;
  wire _2877_;
  wire _2878_;
  wire _2879_;
  wire _2880_;
  wire _2881_;
  wire [63:0] _2882_;
  wire [63:0] _2883_;
  wire [63:0] _2884_;
  wire [63:0] _2885_;
  wire [63:0] _2886_;
  wire [63:0] _2887_;
  wire [63:0] _2888_;
  wire [63:0] _2889_;
  wire [63:0] _2890_;
  wire [63:0] _2891_;
  wire [63:0] _2892_;
  wire [63:0] _2893_;
  wire [8:0] _2894_;
  wire [8:0] _2895_;
  wire [8:0] _2896_;
  wire [8:0] _2897_;
  wire [8:0] _2898_;
  wire [8:0] _2899_;
  wire [8:0] _2900_;
  wire [8:0] _2901_;
  wire [8:0] _2902_;
  wire [8:0] _2903_;
  wire [8:0] _2904_;
  wire [8:0] _2905_;
  wire [8:0] _2906_;
  wire [8:0] _2907_;
  wire [8:0] _2908_;
  wire [8:0] _2909_;
  wire [8:0] _2910_;
  wire [2:0] _2911_;
  wire [2:0] _2912_;
  wire [2:0] _2913_;
  wire [2:0] _2914_;
  wire [2:0] _2915_;
  wire [2:0] _2916_;
  wire [2:0] _2917_;
  wire [2:0] _2918_;
  wire [2:0] _2919_;
  wire [2:0] _2920_;
  wire [2:0] _2921_;
  wire [2:0] _2922_;
  wire [2:0] _2923_;
  wire [2:0] _2924_;
  wire [2:0] _2925_;
  wire [2:0] _2926_;
  wire [2:0] _2927_;
  wire [2:0] _2928_;
  wire [2:0] _2929_;
  wire [2:0] _2930_;
  wire [2:0] _2931_;
  wire [2:0] _2932_;
  wire [2:0] _2933_;
  wire [2:0] _2934_;
  wire [2:0] _2935_;
  wire [2:0] _2936_;
  wire [2:0] _2937_;
  wire [2:0] _2938_;
  wire [2:0] _2939_;
  wire _2940_;
  wire _2941_;
  wire _2942_;
  wire _2943_;
  wire _2944_;
  wire _2945_;
  wire _2946_;
  wire _2947_;
  wire _2948_;
  wire _2949_;
  wire _2950_;
  wire _2951_;
  wire _2952_;
  wire _2953_;
  wire _2954_;
  wire _2955_;
  wire _2956_;
  wire _2957_;
  wire _2958_;
  wire _2959_;
  wire _2960_;
  wire _2961_;
  wire _2962_;
  wire _2963_;
  wire _2964_;
  wire _2965_;
  wire _2966_;
  wire _2967_;
  wire _2968_;
  wire [2:0] _2969_;
  wire [2:0] _2970_;
  wire [2:0] _2971_;
  wire [2:0] _2972_;
  wire [2:0] _2973_;
  wire [2:0] _2974_;
  wire [2:0] _2975_;
  wire [2:0] _2976_;
  wire [2:0] _2977_;
  wire [2:0] _2978_;
  wire [2:0] _2979_;
  wire [2:0] _2980_;
  wire [2:0] _2981_;
  wire [2:0] _2982_;
  wire [2:0] _2983_;
  wire [2:0] _2984_;
  wire [2:0] _2985_;
  wire [2:0] _2986_;
  wire _2987_;
  wire _2988_;
  wire _2989_;
  wire _2990_;
  wire _2991_;
  wire _2992_;
  wire _2993_;
  wire _2994_;
  wire _2995_;
  wire _2996_;
  wire _2997_;
  wire _2998_;
  wire _2999_;
  wire _3000_;
  wire _3001_;
  wire [31:0] _3002_;
  wire _3003_;
  wire _3004_;
  wire _3005_;
  wire [31:0] _3006_;
  wire [2:0] _3007_;
  wire [2:0] _3008_;
  wire [2:0] _3009_;
  wire [5:0] _3010_;
  wire [5:0] _3011_;
  wire [31:0] _3012_;
  wire [1:0] _3013_;
  wire _3014_;
  wire [31:0] _3015_;
  wire [2:0] _3016_;
  wire [1:0] _3017_;
  wire _3018_;
  wire [31:0] _3019_;
  wire _3020_;
  wire [5:0] _3021_;
  wire _3022_;
  wire [31:0] _3023_;
  wire _3024_;
  wire [3:0] _3025_;
  wire [31:0] _3026_;
  wire [31:0] _3027_;
  wire [31:0] _3028_;
  wire _3029_;
  wire [31:0] _3030_;
  wire _3031_;
  wire [2:0] _3032_;
  wire [1:0] _3033_;
  wire _3034_;
  wire [31:0] _3035_;
  wire _3036_;
  wire _3037_;
  wire _3038_;
  wire [5:0] _3039_;
  wire [5:0] _3040_;
  wire [5:0] _3041_;
  wire _3042_;
  wire _3043_;
  wire _3044_;
  wire [31:0] _3045_;
  wire [31:0] _3046_;
  wire [31:0] _3047_;
  wire _3048_;
  wire _3049_;
  wire [1:0] _3050_;
  wire [1:0] _3051_;
  wire [1:0] _3052_;
  wire [3:0] _3053_;
  wire [1:0] _3054_;
  wire [1:0] _3055_;
  wire _3056_;
  wire [1:0] _3057_;
  wire [1:0] _3058_;
  wire _3059_;
  wire [1:0] _3060_;
  wire [1:0] _3061_;
  wire [1:0] _3062_;
  wire [31:0] _3063_;
  wire [31:0] _3064_;
  wire _3065_;
  wire [5:0] _3066_;
  wire [31:0] _3067_;
  wire _3068_;
  wire _3069_;
  wire _3070_;
  wire _3071_;
  wire _3072_;
  wire _3073_;
  wire _3074_;
  wire _3075_;
  wire _3076_;
  wire _3077_;
  wire _3078_;
  wire _3079_;
  wire _3080_;
  wire _3081_;
  wire _3082_;
  wire _3083_;
  wire _3084_;
  wire _3085_;
  wire _3086_;
  wire _3087_;
  wire _3088_;
  wire _3089_;
  wire _3090_;
  wire _3091_;
  wire _3092_;
  wire _3093_;
  wire _3094_;
  wire _3095_;
  wire _3096_;
  wire _3097_;
  wire _3098_;
  wire _3099_;
  wire _3100_;
  wire _3101_;
  wire _3102_;
  wire _3103_;
  wire _3104_;
  wire _3105_;
  wire _3106_;
  wire _3107_;
  wire _3108_;
  wire _3109_;
  wire _3110_;
  wire _3111_;
  wire _3112_;
  wire _3113_;
  wire _3114_;
  wire _3115_;
  wire _3116_;
  wire _3117_;
  wire _3118_;
  wire _3119_;
  wire _3120_;
  wire _3121_;
  wire _3122_;
  wire _3123_;
  wire _3124_;
  wire _3125_;
  wire _3126_;
  wire _3127_;
  wire _3128_;
  wire _3129_;
  wire _3130_;
  wire _3131_;
  wire _3132_;
  wire _3133_;
  wire _3134_;
  wire _3135_;
  wire _3136_;
  wire _3137_;
  wire _3138_;
  wire _3139_;
  wire _3140_;
  wire _3141_;
  wire _3142_;
  wire _3143_;
  wire _3144_;
  wire _3145_;
  wire _3146_;
  wire _3147_;
  wire _3148_;
  wire _3149_;
  wire _3150_;
  wire _3151_;
  wire _3152_;
  wire _3153_;
  wire _3154_;
  wire _3155_;
  wire _3156_;
  wire _3157_;
  wire _3158_;
  wire _3159_;
  wire _3160_;
  wire _3161_;
  wire _3162_;
  wire _3163_;
  wire _3164_;
  wire _3165_;
  wire _3166_;
  wire _3167_;
  wire _3168_;
  wire _3169_;
  wire _3170_;
  wire _3171_;
  wire _3172_;
  wire _3173_;
  wire _3174_;
  wire _3175_;
  wire _3176_;
  wire _3177_;
  wire _3178_;
  wire _3179_;
  wire _3180_;
  wire _3181_;
  wire _3182_;
  wire _3183_;
  wire _3184_;
  wire _3185_;
  wire _3186_;
  wire _3187_;
  wire _3188_;
  wire _3189_;
  wire _3190_;
  wire _3191_;
  wire _3192_;
  wire _3193_;
  wire _3194_;
  wire _3195_;
  wire _3196_;
  wire _3197_;
  wire _3198_;
  wire _3199_;
  wire _3200_;
  wire _3201_;
  wire _3202_;
  wire _3203_;
  wire _3204_;
  wire _3205_;
  wire _3206_;
  wire _3207_;
  wire _3208_;
  wire _3209_;
  wire _3210_;
  wire _3211_;
  wire _3212_;
  wire _3213_;
  wire _3214_;
  wire _3215_;
  wire _3216_;
  wire _3217_;
  wire _3218_;
  wire _3219_;
  wire _3220_;
  wire _3221_;
  wire _3222_;
  wire _3223_;
  wire _3224_;
  wire _3225_;
  wire _3226_;
  wire _3227_;
  wire _3228_;
  wire _3229_;
  wire _3230_;
  wire _3231_;
  wire _3232_;
  wire _3233_;
  wire _3234_;
  wire _3235_;
  wire _3236_;
  wire _3237_;
  wire _3238_;
  wire _3239_;
  wire _3240_;
  wire [31:0] _3241_;
  wire [31:0] _3242_;
  wire _3243_;
  wire _3244_;
  wire _3245_;
  wire _3246_;
  wire _3247_;
  wire _3248_;
  wire _3249_;
  wire _3250_;
  wire _3251_;
  wire _3252_;
  wire _3253_;
  wire _3254_;
  wire _3255_;
  wire _3256_;
  wire _3257_;
  wire _3258_;
  wire _3259_;
  wire _3260_;
  wire _3261_;
  wire _3262_;
  wire _3263_;
  wire _3264_;
  wire _3265_;
  wire _3266_;
  wire _3267_;
  wire _3268_;
  wire _3269_;
  wire _3270_;
  wire [2:0] _3271_;
  wire [2:0] _3272_;
  wire [2:0] _3273_;
  wire [2:0] _3274_;
  wire [2:0] _3275_;
  wire [2:0] _3276_;
  wire [2:0] _3277_;
  wire [2:0] _3278_;
  wire [2:0] _3279_;
  wire [2:0] _3280_;
  wire [2:0] _3281_;
  wire [2:0] _3282_;
  wire [2:0] _3283_;
  wire [2:0] _3284_;
  wire [2:0] _3285_;
  wire [2:0] _3286_;
  wire [2:0] _3287_;
  wire [2:0] _3288_;
  wire [2:0] _3289_;
  wire [2:0] _3290_;
  wire [2:0] _3291_;
  wire [2:0] _3292_;
  wire [2:0] _3293_;
  wire [2:0] _3294_;
  wire [2:0] _3295_;
  wire [2:0] _3296_;
  wire [2:0] _3297_;
  wire [2:0] _3298_;
  wire _3299_;
  wire _3300_;
  wire _3301_;
  wire _3302_;
  wire _3303_;
  wire _3304_;
  wire _3305_;
  wire _3306_;
  wire _3307_;
  wire _3308_;
  wire _3309_;
  wire _3310_;
  wire _3311_;
  wire _3312_;
  wire _3313_;
  wire _3314_;
  wire _3315_;
  wire _3316_;
  wire _3317_;
  wire _3318_;
  wire _3319_;
  wire _3320_;
  wire _3321_;
  wire _3322_;
  wire _3323_;
  wire _3324_;
  wire _3325_;
  wire _3326_;
  wire _3327_;
  wire _3328_;
  wire _3329_;
  wire _3330_;
  wire [2:0] _3331_;
  wire [2:0] _3332_;
  wire [2:0] _3333_;
  wire [2:0] _3334_;
  wire [2:0] _3335_;
  wire [2:0] _3336_;
  wire [2:0] _3337_;
  wire [2:0] _3338_;
  wire [2:0] _3339_;
  wire [2:0] _3340_;
  wire [2:0] _3341_;
  wire [2:0] _3342_;
  wire [2:0] _3343_;
  wire [2:0] _3344_;
  wire [2:0] _3345_;
  wire [2:0] _3346_;
  wire [2:0] _3347_;
  wire [2:0] _3348_;
  wire [2:0] _3349_;
  wire [2:0] _3350_;
  wire [2:0] _3351_;
  wire [2:0] _3352_;
  wire [2:0] _3353_;
  wire [2:0] _3354_;
  wire [2:0] _3355_;
  wire [2:0] _3356_;
  wire [2:0] _3357_;
  wire [2:0] _3358_;
  wire [2:0] _3359_;
  wire [2:0] _3360_;
  wire [2:0] _3361_;
  wire [2:0] _3362_;
  wire [31:0] _3363_;
  wire [31:0] _3364_;
  wire [31:0] _3365_;
  wire [31:0] _3366_;
  wire [31:0] _3367_;
  wire [31:0] _3368_;
  wire [31:0] _3369_;
  wire [31:0] _3370_;
  wire [31:0] _3371_;
  wire [31:0] _3372_;
  wire [31:0] _3373_;
  wire [31:0] _3374_;
  wire [31:0] _3375_;
  wire [31:0] _3376_;
  wire [31:0] _3377_;
  wire [31:0] _3378_;
  wire [31:0] _3379_;
  wire [31:0] _3380_;
  wire [31:0] _3381_;
  wire [31:0] _3382_;
  wire [31:0] _3383_;
  wire _3384_;
  wire _3385_;
  wire _3386_;
  wire _3387_;
  wire _3388_;
  wire _3389_;
  wire _3390_;
  wire _3391_;
  wire _3392_;
  wire _3393_;
  wire _3394_;
  wire _3395_;
  wire _3396_;
  wire _3397_;
  wire _3398_;
  wire _3399_;
  wire _3400_;
  wire _3401_;
  wire _3402_;
  wire _3403_;
  wire _3404_;
  wire _3405_;
  wire _3406_;
  wire _3407_;
  wire _3408_;
  wire _3409_;
  wire _3410_;
  wire _3411_;
  wire _3412_;
  wire _3413_;
  wire _3414_;
  wire _3415_;
  wire _3416_;
  wire _3417_;
  wire _3418_;
  wire _3419_;
  wire _3420_;
  wire _3421_;
  wire _3422_;
  wire _3423_;
  wire _3424_;
  wire _3425_;
  wire _3426_;
  wire _3427_;
  wire _3428_;
  wire _3429_;
  wire _3430_;
  wire _3431_;
  wire _3432_;
  wire _3433_;
  wire _3434_;
  wire _3435_;
  wire _3436_;
  wire _3437_;
  wire _3438_;
  wire _3439_;
  wire _3440_;
  wire _3441_;
  wire _3442_;
  wire _3443_;
  wire _3444_;
  wire _3445_;
  wire _3446_;
  wire _3447_;
  wire _3448_;
  wire _3449_;
  wire _3450_;
  wire _3451_;
  wire _3452_;
  wire _3453_;
  wire _3454_;
  wire _3455_;
  wire _3456_;
  wire _3457_;
  wire _3458_;
  wire _3459_;
  wire _3460_;
  wire _3461_;
  wire _3462_;
  wire _3463_;
  wire _3464_;
  wire _3465_;
  wire _3466_;
  wire _3467_;
  wire _3468_;
  wire _3469_;
  wire _3470_;
  wire _3471_;
  wire _3472_;
  wire _3473_;
  wire _3474_;
  wire _3475_;
  wire _3476_;
  wire _3477_;
  wire _3478_;
  wire _3479_;
  wire _3480_;
  wire _3481_;
  wire _3482_;
  wire _3483_;
  wire _3484_;
  wire _3485_;
  wire [63:0] _3486_;
  wire [63:0] _3487_;
  wire [63:0] _3488_;
  wire [63:0] _3489_;
  wire [63:0] _3490_;
  wire [63:0] _3491_;
  wire [63:0] _3492_;
  wire [63:0] _3493_;
  wire [63:0] _3494_;
  wire [63:0] _3495_;
  wire [63:0] _3496_;
  wire [63:0] _3497_;
  wire [63:0] _3498_;
  wire [63:0] _3499_;
  wire [63:0] _3500_;
  wire [63:0] _3501_;
  wire [63:0] _3502_;
  wire [63:0] _3503_;
  wire [63:0] _3504_;
  wire [63:0] _3505_;
  wire [63:0] _3506_;
  wire [8:0] _3507_;
  wire [8:0] _3508_;
  wire [8:0] _3509_;
  wire [8:0] _3510_;
  wire [8:0] _3511_;
  wire [8:0] _3512_;
  wire [8:0] _3513_;
  wire [8:0] _3514_;
  wire [8:0] _3515_;
  wire [8:0] _3516_;
  wire [8:0] _3517_;
  wire [8:0] _3518_;
  wire [8:0] _3519_;
  wire [8:0] _3520_;
  wire [8:0] _3521_;
  wire [8:0] _3522_;
  wire [8:0] _3523_;
  wire [8:0] _3524_;
  wire [8:0] _3525_;
  wire [8:0] _3526_;
  wire [8:0] _3527_;
  wire [8:0] _3528_;
  wire [8:0] _3529_;
  wire [8:0] _3530_;
  wire [8:0] _3531_;
  wire [8:0] _3532_;
  wire [8:0] _3533_;
  wire [8:0] _3534_;
  wire [8:0] _3535_;
  wire [8:0] _3536_;
  wire [8:0] _3537_;
  wire [8:0] _3538_;
  wire [8:0] _3539_;
  wire [8:0] _3540_;
  wire [2:0] _3541_;
  wire [2:0] _3542_;
  wire [2:0] _3543_;
  wire [2:0] _3544_;
  wire [2:0] _3545_;
  wire [2:0] _3546_;
  wire [2:0] _3547_;
  wire [2:0] _3548_;
  wire [2:0] _3549_;
  wire [2:0] _3550_;
  wire [2:0] _3551_;
  wire [2:0] _3552_;
  wire [2:0] _3553_;
  wire [2:0] _3554_;
  wire [2:0] _3555_;
  wire [2:0] _3556_;
  wire [2:0] _3557_;
  wire [2:0] _3558_;
  wire [2:0] _3559_;
  wire [2:0] _3560_;
  wire [2:0] _3561_;
  wire [2:0] _3562_;
  wire [2:0] _3563_;
  wire [2:0] _3564_;
  wire [2:0] _3565_;
  wire [2:0] _3566_;
  wire [2:0] _3567_;
  wire [2:0] _3568_;
  wire [2:0] _3569_;
  wire [2:0] _3570_;
  wire [2:0] _3571_;
  wire [2:0] _3572_;
  wire [2:0] _3573_;
  wire [2:0] _3574_;
  wire [2:0] _3575_;
  wire [2:0] _3576_;
  wire [2:0] _3577_;
  wire [2:0] _3578_;
  wire [2:0] _3579_;
  wire [2:0] _3580_;
  wire [2:0] _3581_;
  wire [2:0] _3582_;
  wire [2:0] _3583_;
  wire [2:0] _3584_;
  wire [2:0] _3585_;
  wire [2:0] _3586_;
  wire [2:0] _3587_;
  wire [2:0] _3588_;
  wire [2:0] _3589_;
  wire [2:0] _3590_;
  wire [2:0] _3591_;
  wire [2:0] _3592_;
  wire [2:0] _3593_;
  wire [2:0] _3594_;
  wire [2:0] _3595_;
  wire [2:0] _3596_;
  wire [2:0] _3597_;
  wire [2:0] _3598_;
  wire _3599_;
  wire _3600_;
  wire _3601_;
  wire _3602_;
  wire _3603_;
  wire _3604_;
  wire _3605_;
  wire _3606_;
  wire _3607_;
  wire _3608_;
  wire _3609_;
  wire _3610_;
  wire _3611_;
  wire _3612_;
  wire _3613_;
  wire _3614_;
  wire _3615_;
  wire _3616_;
  wire _3617_;
  wire _3618_;
  wire _3619_;
  wire _3620_;
  wire _3621_;
  wire _3622_;
  wire _3623_;
  wire _3624_;
  wire _3625_;
  wire _3626_;
  wire _3627_;
  wire _3628_;
  wire _3629_;
  wire _3630_;
  wire _3631_;
  wire _3632_;
  wire _3633_;
  wire _3634_;
  wire _3635_;
  wire _3636_;
  wire _3637_;
  wire _3638_;
  wire _3639_;
  wire _3640_;
  wire _3641_;
  wire _3642_;
  wire _3643_;
  wire _3644_;
  wire _3645_;
  wire _3646_;
  wire _3647_;
  wire _3648_;
  wire _3649_;
  wire _3650_;
  wire _3651_;
  wire _3652_;
  wire _3653_;
  wire _3654_;
  wire _3655_;
  wire _3656_;
  wire _3657_;
  wire _3658_;
  wire _3659_;
  wire _3660_;
  wire [2:0] _3661_;
  wire [2:0] _3662_;
  wire [2:0] _3663_;
  wire [2:0] _3664_;
  wire [2:0] _3665_;
  wire [2:0] _3666_;
  wire [2:0] _3667_;
  wire [2:0] _3668_;
  wire [2:0] _3669_;
  wire [2:0] _3670_;
  wire [2:0] _3671_;
  wire [2:0] _3672_;
  wire [2:0] _3673_;
  wire [2:0] _3674_;
  wire [2:0] _3675_;
  wire [2:0] _3676_;
  wire [2:0] _3677_;
  wire [2:0] _3678_;
  wire [2:0] _3679_;
  wire [2:0] _3680_;
  wire [2:0] _3681_;
  wire [2:0] _3682_;
  wire [2:0] _3683_;
  wire [2:0] _3684_;
  wire [2:0] _3685_;
  wire [2:0] _3686_;
  wire [2:0] _3687_;
  wire [2:0] _3688_;
  wire [2:0] _3689_;
  wire [2:0] _3690_;
  wire [2:0] _3691_;
  wire [2:0] _3692_;
  wire [2:0] _3693_;
  wire [2:0] _3694_;
  wire [2:0] _3695_;
  wire [2:0] _3696_;
  wire _3697_;
  wire _3698_;
  wire _3699_;
  wire _3700_;
  wire _3701_;
  wire _3702_;
  wire _3703_;
  wire _3704_;
  wire _3705_;
  wire _3706_;
  wire _3707_;
  wire _3708_;
  wire _3709_;
  wire _3710_;
  wire _3711_;
  wire _3712_;
  wire _3713_;
  wire _3714_;
  wire _3715_;
  wire _3716_;
  wire _3717_;
  wire _3718_;
  wire _3719_;
  wire _3720_;
  wire _3721_;
  wire _3722_;
  wire _3723_;
  wire _3724_;
  wire _3725_;
  wire _3726_;
  wire _3727_;
  wire [31:0] _3728_;
  wire _3729_;
  wire _3730_;
  wire _3731_;
  wire _3732_;
  wire _3733_;
  wire _3734_;
  wire _3735_;
  wire _3736_;
  wire _3737_;
  wire _3738_;
  wire _3739_;
  wire _3740_;
  wire _3741_;
  wire _3742_;
  wire _3743_;
  wire _3744_;
  wire _3745_;
  wire _3746_;
  wire _3747_;
  wire _3748_;
  wire _3749_;
  wire _3750_;
  wire _3751_;
  wire _3752_;
  wire _3753_;
  wire _3754_;
  wire _3755_;
  wire _3756_;
  wire _3757_;
  wire _3758_;
  wire _3759_;
  wire [31:0] _3760_;
  wire [31:0] _3761_;
  wire [31:0] _3762_;
  wire _3763_;
  wire _3764_;
  wire _3765_;
  wire _3766_;
  wire _3767_;
  wire _3768_;
  wire _3769_;
  wire _3770_;
  wire _3771_;
  wire _3772_;
  wire _3773_;
  wire _3774_;
  wire [31:0] _3775_;
  wire _3776_;
  wire _3777_;
  wire _3778_;
  wire _3779_;
  wire [31:0] _3780_;
  wire [31:0] _3781_;
  wire _3782_;
  wire _3783_;
  wire _3784_;
  wire _3785_;
  wire _3786_;
  wire _3787_;
  wire _3788_;
  wire _3789_;
  wire [2:0] _3790_;
  wire [2:0] _3791_;
  wire [2:0] _3792_;
  wire [2:0] _3793_;
  wire [31:0] _3794_;
  wire [31:0] _3795_;
  wire [31:0] _3796_;
  wire [31:0] _3797_;
  wire _3798_;
  wire _3799_;
  wire _3800_;
  wire _3801_;
  wire [5:0] _3802_;
  wire [5:0] _3803_;
  wire [5:0] _3804_;
  wire [5:0] _3805_;
  wire _3806_;
  wire _3807_;
  wire _3808_;
  wire _3809_;
  wire [31:0] _3810_;
  wire [31:0] _3811_;
  wire [31:0] _3812_;
  wire [31:0] _3813_;
  wire _3814_;
  wire _3815_;
  wire _3816_;
  wire _3817_;
  wire [1:0] _3818_;
  wire [1:0] _3819_;
  wire [1:0] _3820_;
  wire [1:0] _3821_;
  wire _3822_;
  wire _3823_;
  wire [30:0] _3824_;
  wire [30:0] _3825_;
  wire _3826_;
  wire _3827_;
  wire [30:0] _3828_;
  wire [30:0] _3829_;
  wire _3830_;
  wire _3831_;
  wire _3832_;
  wire _3833_;
  wire _3834_;
  wire _3835_;
  wire _3836_;
  wire _3837_;
  wire _3838_;
  wire _3839_;
  wire _3840_;
  wire _3841_;
  wire _3842_;
  wire _3843_;
  wire [28:0] _3844_;
  wire [28:0] _3845_;
  wire _3846_;
  wire _3847_;
  wire _3848_;
  wire _3849_;
  wire _3850_;
  wire _3851_;
  wire _3852_;
  wire _3853_;
  wire _3854_;
  wire _3855_;
  wire _3856_;
  wire _3857_;
  wire _3858_;
  wire _3859_;
  wire _3860_;
  wire _3861_;
  wire _3862_;
  wire _3863_;
  wire _3864_;
  wire _3865_;
  wire _3866_;
  wire _3867_;
  wire _3868_;
  wire _3869_;
  wire _3870_;
  wire _3871_;
  wire _3872_;
  wire _3873_;
  wire _3874_;
  wire _3875_;
  wire _3876_;
  wire _3877_;
  wire _3878_;
  wire _3879_;
  wire _3880_;
  wire _3881_;
  wire _3882_;
  wire _3883_;
  wire _3884_;
  wire _3885_;
  wire _3886_;
  wire _3887_;
  wire _3888_;
  wire _3889_;
  wire _3890_;
  wire _3891_;
  wire _3892_;
  wire _3893_;
  wire _3894_;
  wire _3895_;
  wire _3896_;
  wire _3897_;
  wire _3898_;
  wire _3899_;
  wire _3900_;
  wire _3901_;
  wire _3902_;
  wire _3903_;
  wire _3904_;
  wire _3905_;
  wire _3906_;
  wire _3907_;
  wire _3908_;
  wire _3909_;
  wire _3910_;
  wire _3911_;
  wire _3912_;
  wire _3913_;
  wire _3914_;
  wire _3915_;
  wire _3916_;
  wire _3917_;
  wire _3918_;
  wire _3919_;
  wire _3920_;
  wire _3921_;
  wire _3922_;
  wire _3923_;
  wire _3924_;
  wire _3925_;
  wire _3926_;
  wire _3927_;
  wire _3928_;
  wire _3929_;
  wire _3930_;
  wire _3931_;
  wire _3932_;
  wire _3933_;
  wire _3934_;
  wire _3935_;
  wire _3936_;
  wire _3937_;
  wire _3938_;
  wire _3939_;
  wire _3940_;
  wire _3941_;
  wire _3942_;
  wire _3943_;
  wire _3944_;
  wire _3945_;
  wire _3946_;
  wire _3947_;
  wire _3948_;
  wire _3949_;
  wire _3950_;
  wire _3951_;
  wire _3952_;
  wire _3953_;
  wire _3954_;
  wire _3955_;
  wire _3956_;
  wire _3957_;
  wire _3958_;
  wire _3959_;
  wire _3960_;
  wire _3961_;
  wire _3962_;
  wire _3963_;
  wire _3964_;
  wire _3965_;
  wire [31:0] _3966_;
  input [31:0] boot_addr_i;
  wire [31:0] boot_addr_i;
  input [31:0] boot_addr_i_t0;
  wire [31:0] boot_addr_i_t0;
  input branch_i;
  wire branch_i;
  input branch_i_t0;
  wire branch_i_t0;
  input branch_taken_i;
  wire branch_taken_i;
  input branch_taken_i_t0;
  wire branch_taken_i_t0;
  input clk_i;
  wire clk_i;
  wire cpuctrl_err;
  wire cpuctrl_err_t0;
  wire [5:0] cpuctrl_q;
  wire [5:0] cpuctrl_q_t0;
  wire cpuctrl_we;
  wire cpuctrl_we_t0;
  input csr_access_i;
  wire csr_access_i;
  input csr_access_i_t0;
  wire csr_access_i_t0;
  input [11:0] csr_addr_i;
  wire [11:0] csr_addr_i;
  input [11:0] csr_addr_i_t0;
  wire [11:0] csr_addr_i_t0;
  output [31:0] csr_depc_o;
  wire [31:0] csr_depc_o;
  output [31:0] csr_depc_o_t0;
  wire [31:0] csr_depc_o_t0;
  input [5:0] csr_mcause_i;
  wire [5:0] csr_mcause_i;
  input [5:0] csr_mcause_i_t0;
  wire [5:0] csr_mcause_i_t0;
  output [31:0] csr_mepc_o;
  wire [31:0] csr_mepc_o;
  output [31:0] csr_mepc_o_t0;
  wire [31:0] csr_mepc_o_t0;
  output csr_mstatus_mie_o;
  wire csr_mstatus_mie_o;
  output csr_mstatus_mie_o_t0;
  wire csr_mstatus_mie_o_t0;
  output csr_mstatus_tw_o;
  wire csr_mstatus_tw_o;
  output csr_mstatus_tw_o_t0;
  wire csr_mstatus_tw_o_t0;
  input [31:0] csr_mtval_i;
  wire [31:0] csr_mtval_i;
  input [31:0] csr_mtval_i_t0;
  wire [31:0] csr_mtval_i_t0;
  input csr_mtvec_init_i;
  wire csr_mtvec_init_i;
  input csr_mtvec_init_i_t0;
  wire csr_mtvec_init_i_t0;
  output [31:0] csr_mtvec_o;
  wire [31:0] csr_mtvec_o;
  output [31:0] csr_mtvec_o_t0;
  wire [31:0] csr_mtvec_o_t0;
  input csr_op_en_i;
  wire csr_op_en_i;
  input csr_op_en_i_t0;
  wire csr_op_en_i_t0;
  input [1:0] csr_op_i;
  wire [1:0] csr_op_i;
  input [1:0] csr_op_i_t0;
  wire [1:0] csr_op_i_t0;
  output [135:0] csr_pmp_addr_o;
  wire [135:0] csr_pmp_addr_o;
  output [135:0] csr_pmp_addr_o_t0;
  wire [135:0] csr_pmp_addr_o_t0;
  output [23:0] csr_pmp_cfg_o;
  wire [23:0] csr_pmp_cfg_o;
  output [23:0] csr_pmp_cfg_o_t0;
  wire [23:0] csr_pmp_cfg_o_t0;
  output [2:0] csr_pmp_mseccfg_o;
  wire [2:0] csr_pmp_mseccfg_o;
  output [2:0] csr_pmp_mseccfg_o_t0;
  wire [2:0] csr_pmp_mseccfg_o_t0;
  output [31:0] csr_rdata_o;
  wire [31:0] csr_rdata_o;
  output [31:0] csr_rdata_o_t0;
  wire [31:0] csr_rdata_o_t0;
  input csr_restore_dret_i;
  wire csr_restore_dret_i;
  input csr_restore_dret_i_t0;
  wire csr_restore_dret_i_t0;
  input csr_restore_mret_i;
  wire csr_restore_mret_i;
  input csr_restore_mret_i_t0;
  wire csr_restore_mret_i_t0;
  input csr_save_cause_i;
  wire csr_save_cause_i;
  input csr_save_cause_i_t0;
  wire csr_save_cause_i_t0;
  input csr_save_id_i;
  wire csr_save_id_i;
  input csr_save_id_i_t0;
  wire csr_save_id_i_t0;
  input csr_save_if_i;
  wire csr_save_if_i;
  input csr_save_if_i_t0;
  wire csr_save_if_i_t0;
  input csr_save_wb_i;
  wire csr_save_wb_i;
  input csr_save_wb_i_t0;
  wire csr_save_wb_i_t0;
  output csr_shadow_err_o;
  wire csr_shadow_err_o;
  output csr_shadow_err_o_t0;
  wire csr_shadow_err_o_t0;
  input [31:0] csr_wdata_i;
  wire [31:0] csr_wdata_i;
  input [31:0] csr_wdata_i_t0;
  wire [31:0] csr_wdata_i_t0;
  wire [31:0] csr_wdata_int;
  wire [31:0] csr_wdata_int_t0;
  wire csr_we_int;
  wire csr_we_int_t0;
  wire csr_wr;
  wire csr_wr_t0;
  output data_ind_timing_o;
  wire data_ind_timing_o;
  output data_ind_timing_o_t0;
  wire data_ind_timing_o_t0;
  wire [31:0] dcsr_d;
  wire [31:0] dcsr_d_t0;
  wire dcsr_en;
  wire dcsr_en_t0;
  wire [31:0] dcsr_q;
  wire [31:0] dcsr_q_t0;
  input [2:0] debug_cause_i;
  wire [2:0] debug_cause_i;
  input [2:0] debug_cause_i_t0;
  wire [2:0] debug_cause_i_t0;
  input debug_csr_save_i;
  wire debug_csr_save_i;
  input debug_csr_save_i_t0;
  wire debug_csr_save_i_t0;
  output debug_ebreakm_o;
  wire debug_ebreakm_o;
  output debug_ebreakm_o_t0;
  wire debug_ebreakm_o_t0;
  output debug_ebreaku_o;
  wire debug_ebreaku_o;
  output debug_ebreaku_o_t0;
  wire debug_ebreaku_o_t0;
  input debug_mode_i;
  wire debug_mode_i;
  input debug_mode_i_t0;
  wire debug_mode_i_t0;
  output debug_single_step_o;
  wire debug_single_step_o;
  output debug_single_step_o_t0;
  wire debug_single_step_o_t0;
  wire [31:0] depc_d;
  wire [31:0] depc_d_t0;
  wire depc_en;
  wire depc_en_t0;
  input div_wait_i;
  wire div_wait_i;
  input div_wait_i_t0;
  wire div_wait_i_t0;
  wire dscratch0_en;
  wire dscratch0_en_t0;
  wire [31:0] dscratch0_q;
  wire [31:0] dscratch0_q_t0;
  wire dscratch1_en;
  wire dscratch1_en_t0;
  wire [31:0] dscratch1_q;
  wire [31:0] dscratch1_q_t0;
  input dside_wait_i;
  wire dside_wait_i;
  input dside_wait_i_t0;
  wire dside_wait_i_t0;
  output dummy_instr_en_o;
  wire dummy_instr_en_o;
  output dummy_instr_en_o_t0;
  wire dummy_instr_en_o_t0;
  output [2:0] dummy_instr_mask_o;
  wire [2:0] dummy_instr_mask_o;
  output [2:0] dummy_instr_mask_o_t0;
  wire [2:0] dummy_instr_mask_o_t0;
  output dummy_instr_seed_en_o;
  wire dummy_instr_seed_en_o;
  output dummy_instr_seed_en_o_t0;
  wire dummy_instr_seed_en_o_t0;
  output [31:0] dummy_instr_seed_o;
  wire [31:0] dummy_instr_seed_o;
  output [31:0] dummy_instr_seed_o_t0;
  wire [31:0] dummy_instr_seed_o_t0;
  wire \gen_trigger_regs.selected_tmatch_control ;
  wire \gen_trigger_regs.selected_tmatch_control_t0 ;
  wire [31:0] \gen_trigger_regs.selected_tmatch_value ;
  wire [31:0] \gen_trigger_regs.selected_tmatch_value_t0 ;
  wire \gen_trigger_regs.tmatch_control_we ;
  wire \gen_trigger_regs.tmatch_control_we_t0 ;
  wire \gen_trigger_regs.tmatch_value_we ;
  wire \gen_trigger_regs.tmatch_value_we_t0 ;
  wire \gen_trigger_regs.tselect_d ;
  wire \gen_trigger_regs.tselect_d_t0 ;
  wire \gen_trigger_regs.tselect_q ;
  wire \gen_trigger_regs.tselect_q_t0 ;
  wire \gen_trigger_regs.tselect_we ;
  wire \gen_trigger_regs.tselect_we_t0 ;
  input [31:0] hart_id_i;
  wire [31:0] hart_id_i;
  input [31:0] hart_id_i_t0;
  wire [31:0] hart_id_i_t0;
  output icache_enable_o;
  wire icache_enable_o;
  output icache_enable_o_t0;
  wire icache_enable_o_t0;
  wire illegal_csr;
  output illegal_csr_insn_o;
  wire illegal_csr_insn_o;
  output illegal_csr_insn_o_t0;
  wire illegal_csr_insn_o_t0;
  wire illegal_csr_priv;
  wire illegal_csr_priv_t0;
  wire illegal_csr_t0;
  wire illegal_csr_write;
  wire illegal_csr_write_t0;
  input instr_ret_compressed_i;
  wire instr_ret_compressed_i;
  input instr_ret_compressed_i_t0;
  wire instr_ret_compressed_i_t0;
  input instr_ret_i;
  wire instr_ret_i;
  input instr_ret_i_t0;
  wire instr_ret_i_t0;
  input irq_external_i;
  wire irq_external_i;
  input irq_external_i_t0;
  wire irq_external_i_t0;
  input [14:0] irq_fast_i;
  wire [14:0] irq_fast_i;
  input [14:0] irq_fast_i_t0;
  wire [14:0] irq_fast_i_t0;
  output irq_pending_o;
  wire irq_pending_o;
  output irq_pending_o_t0;
  wire irq_pending_o_t0;
  input irq_software_i;
  wire irq_software_i;
  input irq_software_i_t0;
  wire irq_software_i_t0;
  input irq_timer_i;
  wire irq_timer_i;
  input irq_timer_i_t0;
  wire irq_timer_i_t0;
  output [17:0] irqs_o;
  wire [17:0] irqs_o;
  output [17:0] irqs_o_t0;
  wire [17:0] irqs_o_t0;
  input iside_wait_i;
  wire iside_wait_i;
  input iside_wait_i_t0;
  wire iside_wait_i_t0;
  input jump_i;
  wire jump_i;
  input jump_i_t0;
  wire jump_i_t0;
  wire [5:0] mcause_d;
  wire [5:0] mcause_d_t0;
  wire mcause_en;
  wire mcause_en_t0;
  wire [5:0] mcause_q;
  wire [5:0] mcause_q_t0;
  wire [31:0] mcountinhibit;
  wire [31:0] mcountinhibit_t0;
  wire mcountinhibit_we;
  wire mcountinhibit_we_t0;
  input mem_load_i;
  wire mem_load_i;
  input mem_load_i_t0;
  wire mem_load_i_t0;
  input mem_store_i;
  wire mem_store_i;
  input mem_store_i_t0;
  wire mem_store_i_t0;
  wire [31:0] mepc_d;
  wire [31:0] mepc_d_t0;
  wire mepc_en;
  wire mepc_en_t0;
  wire [63:0] \mhpmcounter[0] ;
  wire [63:0] \mhpmcounter[0]_t0 ;
  wire [63:0] \mhpmcounter[10] ;
  wire [63:0] \mhpmcounter[10]_t0 ;
  wire [63:0] \mhpmcounter[11] ;
  wire [63:0] \mhpmcounter[11]_t0 ;
  wire [63:0] \mhpmcounter[12] ;
  wire [63:0] \mhpmcounter[12]_t0 ;
  wire [63:0] \mhpmcounter[2] ;
  wire [63:0] \mhpmcounter[2]_t0 ;
  wire [63:0] \mhpmcounter[3] ;
  wire [63:0] \mhpmcounter[3]_t0 ;
  wire [63:0] \mhpmcounter[4] ;
  wire [63:0] \mhpmcounter[4]_t0 ;
  wire [63:0] \mhpmcounter[5] ;
  wire [63:0] \mhpmcounter[5]_t0 ;
  wire [63:0] \mhpmcounter[6] ;
  wire [63:0] \mhpmcounter[6]_t0 ;
  wire [63:0] \mhpmcounter[7] ;
  wire [63:0] \mhpmcounter[7]_t0 ;
  wire [63:0] \mhpmcounter[8] ;
  wire [63:0] \mhpmcounter[8]_t0 ;
  wire [63:0] \mhpmcounter[9] ;
  wire [63:0] \mhpmcounter[9]_t0 ;
  wire [31:0] mhpmcounter_we;
  wire [31:0] mhpmcounter_we_t0;
  wire [31:0] mhpmcounterh_we;
  wire [31:0] mhpmcounterh_we_t0;
  wire mie_en;
  wire mie_en_t0;
  wire [17:0] mie_q;
  wire [17:0] mie_q_t0;
  wire mscratch_en;
  wire mscratch_en_t0;
  wire [31:0] mscratch_q;
  wire [31:0] mscratch_q_t0;
  wire [5:0] mstack_cause_q;
  wire [5:0] mstack_cause_q_t0;
  wire mstack_en;
  wire mstack_en_t0;
  wire [31:0] mstack_epc_q;
  wire [31:0] mstack_epc_q_t0;
  wire [2:0] mstack_q;
  wire [2:0] mstack_q_t0;
  wire [5:0] mstatus_d;
  wire [5:0] mstatus_d_t0;
  wire mstatus_en;
  wire mstatus_en_t0;
  wire mstatus_err;
  wire mstatus_err_t0;
  wire [5:0] mstatus_q;
  wire [5:0] mstatus_q_t0;
  wire [31:0] mtval_d;
  wire [31:0] mtval_d_t0;
  wire mtval_en;
  wire mtval_en_t0;
  wire [31:0] mtval_q;
  wire [31:0] mtval_q_t0;
  wire [31:0] mtvec_d;
  wire [31:0] mtvec_d_t0;
  wire mtvec_en;
  wire mtvec_en_t0;
  wire mtvec_err;
  wire mtvec_err_t0;
  input mul_wait_i;
  wire mul_wait_i;
  input mul_wait_i_t0;
  wire mul_wait_i_t0;
  input nmi_mode_i;
  wire nmi_mode_i;
  input nmi_mode_i_t0;
  wire nmi_mode_i_t0;
  input [31:0] pc_id_i;
  wire [31:0] pc_id_i;
  input [31:0] pc_id_i_t0;
  wire [31:0] pc_id_i_t0;
  input [31:0] pc_if_i;
  wire [31:0] pc_if_i;
  input [31:0] pc_if_i_t0;
  wire [31:0] pc_if_i_t0;
  input [31:0] pc_wb_i;
  wire [31:0] pc_wb_i;
  input [31:0] pc_wb_i_t0;
  wire [31:0] pc_wb_i_t0;
  output [1:0] priv_mode_id_o;
  reg [1:0] priv_mode_id_o;
  output [1:0] priv_mode_id_o_t0;
  reg [1:0] priv_mode_id_o_t0;
  output [1:0] priv_mode_if_o;
  wire [1:0] priv_mode_if_o;
  output [1:0] priv_mode_if_o_t0;
  wire [1:0] priv_mode_if_o_t0;
  output [1:0] priv_mode_lsu_o;
  wire [1:0] priv_mode_lsu_o;
  output [1:0] priv_mode_lsu_o_t0;
  wire [1:0] priv_mode_lsu_o_t0;
  input rst_ni;
  wire rst_ni;
  output trigger_match_o;
  wire trigger_match_o;
  output trigger_match_o_t0;
  wire trigger_match_o_t0;
  assign illegal_csr_insn_o = csr_access_i & _3778_;
  assign _0117_ = _0353_ & csr_rdata_o;
  assign _0119_ = csr_wr & csr_op_en_i;
  assign csr_we_int = _0119_ & _3763_;
  assign irqs_o = { irq_software_i, irq_timer_i, irq_external_i, irq_fast_i } & mie_q;
  assign _0122_ = instr_ret_i & _3764_;
  assign _0124_ = dside_wait_i & _3765_;
  assign _0126_ = iside_wait_i & _3766_;
  assign _0128_ = mem_load_i & _3767_;
  assign _0130_ = mem_store_i & _3768_;
  assign _0132_ = jump_i & _3769_;
  assign _0134_ = branch_i & _3770_;
  assign _0136_ = branch_taken_i & _3771_;
  assign _0138_ = instr_ret_compressed_i & _3772_;
  assign _0140_ = mul_wait_i & _3773_;
  assign _0142_ = div_wait_i & _3774_;
  assign _0144_ = csr_we_int & debug_mode_i;
  assign \gen_trigger_regs.tselect_we  = _0144_ & _3737_;
  assign \gen_trigger_regs.tmatch_control_we  = _0148_ & _3740_;
  assign _0146_ = _3739_ & csr_we_int;
  assign _0148_ = _0146_ & debug_mode_i;
  assign \gen_trigger_regs.tmatch_value_we  = _0148_ & _3742_;
  assign trigger_match_o = \gen_trigger_regs.selected_tmatch_control  & _3744_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) priv_mode_id_o_t0 <= 2'h0;
    else priv_mode_id_o_t0 <= priv_mode_if_o_t0;
  assign _0164_ = ~ mcountinhibit_we;
  assign _2764_ = { csr_wdata_int[12:2], csr_wdata_int[0] } ^ { mcountinhibit[12:2], mcountinhibit[0] };
  assign _2049_ = { csr_wdata_int_t0[12:2], csr_wdata_int_t0[0] } | { mcountinhibit_t0[12:2], mcountinhibit_t0[0] };
  assign _2050_ = _2764_ | _2049_;
  assign _0641_ = { mcountinhibit_we, mcountinhibit_we, mcountinhibit_we, mcountinhibit_we, mcountinhibit_we, mcountinhibit_we, mcountinhibit_we, mcountinhibit_we, mcountinhibit_we, mcountinhibit_we, mcountinhibit_we, mcountinhibit_we } & { csr_wdata_int_t0[12:2], csr_wdata_int_t0[0] };
  assign _0642_ = { _0164_, _0164_, _0164_, _0164_, _0164_, _0164_, _0164_, _0164_, _0164_, _0164_, _0164_, _0164_ } & { mcountinhibit_t0[12:2], mcountinhibit_t0[0] };
  assign _0643_ = _2050_ & { mcountinhibit_we_t0, mcountinhibit_we_t0, mcountinhibit_we_t0, mcountinhibit_we_t0, mcountinhibit_we_t0, mcountinhibit_we_t0, mcountinhibit_we_t0, mcountinhibit_we_t0, mcountinhibit_we_t0, mcountinhibit_we_t0, mcountinhibit_we_t0, mcountinhibit_we_t0 };
  assign _2051_ = _0641_ | _0642_;
  assign _2052_ = _2051_ | _0643_;
  reg [11:0] _4000_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) _4000_ <= 12'h000;
    else _4000_ <= _2052_;
  assign { mcountinhibit_t0[12:2], mcountinhibit_t0[0] } = _4000_;
  assign _0115_ = 32'd0 & _0348_;
  assign _0572_ = csr_access_i_t0 & _3778_;
  assign _0575_ = csr_wdata_i_t0 & csr_rdata_o;
  assign _0578_ = csr_wr_t0 & csr_op_en_i;
  assign _0581_ = _0120_ & _3763_;
  assign _0584_ = { irq_software_i_t0, irq_timer_i_t0, irq_external_i_t0, irq_fast_i_t0 } & mie_q;
  assign _0587_ = instr_ret_i_t0 & _3764_;
  assign _0590_ = dside_wait_i_t0 & _3765_;
  assign _0593_ = iside_wait_i_t0 & _3766_;
  assign _0596_ = mem_load_i_t0 & _3767_;
  assign _0599_ = mem_store_i_t0 & _3768_;
  assign _0602_ = jump_i_t0 & _3769_;
  assign _0605_ = branch_i_t0 & _3770_;
  assign _0608_ = branch_taken_i_t0 & _3771_;
  assign _0611_ = instr_ret_compressed_i_t0 & _3772_;
  assign _0614_ = mul_wait_i_t0 & _3773_;
  assign _0617_ = div_wait_i_t0 & _3774_;
  assign _0620_ = csr_we_int_t0 & debug_mode_i;
  assign _0623_ = _0145_ & _3737_;
  assign _0626_ = _0149_ & _3740_;
  assign _0629_ = \gen_trigger_regs.tselect_q_t0  & csr_we_int;
  assign _0632_ = _0147_ & debug_mode_i;
  assign _0635_ = _0149_ & _3742_;
  assign _0638_ = \gen_trigger_regs.selected_tmatch_control_t0  & _3744_;
  assign _0573_ = _3779_ & csr_access_i;
  assign _0579_ = csr_op_en_i_t0 & csr_wr;
  assign _0582_ = illegal_csr_insn_o_t0 & _0119_;
  assign _0585_ = mie_q_t0 & { irq_software_i, irq_timer_i, irq_external_i, irq_fast_i };
  assign _0588_ = mcountinhibit_t0[2] & instr_ret_i;
  assign _0591_ = mcountinhibit_t0[3] & dside_wait_i;
  assign _0594_ = mcountinhibit_t0[4] & iside_wait_i;
  assign _0597_ = mcountinhibit_t0[5] & mem_load_i;
  assign _0600_ = mcountinhibit_t0[6] & mem_store_i;
  assign _0603_ = mcountinhibit_t0[7] & jump_i;
  assign _0606_ = mcountinhibit_t0[8] & branch_i;
  assign _0609_ = mcountinhibit_t0[9] & branch_taken_i;
  assign _0612_ = mcountinhibit_t0[10] & instr_ret_compressed_i;
  assign _0615_ = mcountinhibit_t0[11] & mul_wait_i;
  assign _0618_ = mcountinhibit_t0[12] & div_wait_i;
  assign _0621_ = debug_mode_i_t0 & csr_we_int;
  assign _0624_ = _3738_ & _0144_;
  assign _0627_ = _3741_ & _0148_;
  assign _0630_ = csr_we_int_t0 & _3739_;
  assign _0633_ = debug_mode_i_t0 & _0146_;
  assign _0636_ = _3743_ & _0148_;
  assign _0639_ = _3745_ & \gen_trigger_regs.selected_tmatch_control ;
  assign _0571_ = 32'd0 & _3762_;
  assign _0574_ = csr_access_i_t0 & _3779_;
  assign _0580_ = csr_wr_t0 & csr_op_en_i_t0;
  assign _0583_ = _0120_ & illegal_csr_insn_o_t0;
  assign _0586_ = { irq_software_i_t0, irq_timer_i_t0, irq_external_i_t0, irq_fast_i_t0 } & mie_q_t0;
  assign _0589_ = instr_ret_i_t0 & mcountinhibit_t0[2];
  assign _0592_ = dside_wait_i_t0 & mcountinhibit_t0[3];
  assign _0595_ = iside_wait_i_t0 & mcountinhibit_t0[4];
  assign _0598_ = mem_load_i_t0 & mcountinhibit_t0[5];
  assign _0601_ = mem_store_i_t0 & mcountinhibit_t0[6];
  assign _0604_ = jump_i_t0 & mcountinhibit_t0[7];
  assign _0607_ = branch_i_t0 & mcountinhibit_t0[8];
  assign _0610_ = branch_taken_i_t0 & mcountinhibit_t0[9];
  assign _0613_ = instr_ret_compressed_i_t0 & mcountinhibit_t0[10];
  assign _0616_ = mul_wait_i_t0 & mcountinhibit_t0[11];
  assign _0619_ = div_wait_i_t0 & mcountinhibit_t0[12];
  assign _0622_ = csr_we_int_t0 & debug_mode_i_t0;
  assign _0625_ = _0145_ & _3738_;
  assign _0628_ = _0149_ & _3741_;
  assign _0631_ = \gen_trigger_regs.tselect_q_t0  & csr_we_int_t0;
  assign _0634_ = _0147_ & debug_mode_i_t0;
  assign _0637_ = _0149_ & _3743_;
  assign _0640_ = \gen_trigger_regs.selected_tmatch_control_t0  & _3745_;
  assign _2025_ = _0115_ | _0571_;
  assign _2026_ = _0572_ | _0573_;
  assign _2027_ = _0575_ | _0576_;
  assign _2028_ = _0578_ | _0579_;
  assign _2029_ = _0581_ | _0582_;
  assign _2030_ = _0584_ | _0585_;
  assign _2031_ = _0587_ | _0588_;
  assign _2032_ = _0590_ | _0591_;
  assign _2033_ = _0593_ | _0594_;
  assign _2034_ = _0596_ | _0597_;
  assign _2035_ = _0599_ | _0600_;
  assign _2036_ = _0602_ | _0603_;
  assign _2037_ = _0605_ | _0606_;
  assign _2038_ = _0608_ | _0609_;
  assign _2039_ = _0611_ | _0612_;
  assign _2040_ = _0614_ | _0615_;
  assign _2041_ = _0617_ | _0618_;
  assign _2042_ = _0620_ | _0621_;
  assign _2043_ = _0623_ | _0624_;
  assign _2044_ = _0626_ | _0627_;
  assign _2045_ = _0629_ | _0630_;
  assign _2046_ = _0632_ | _0633_;
  assign _2047_ = _0635_ | _0636_;
  assign _2048_ = _0638_ | _0639_;
  assign _0116_ = _2025_ | _0571_;
  assign illegal_csr_insn_o_t0 = _2026_ | _0574_;
  assign _0118_ = _2027_ | _0577_;
  assign _0120_ = _2028_ | _0580_;
  assign csr_we_int_t0 = _2029_ | _0583_;
  assign irqs_o_t0 = _2030_ | _0586_;
  assign _0123_ = _2031_ | _0589_;
  assign _0125_ = _2032_ | _0592_;
  assign _0127_ = _2033_ | _0595_;
  assign _0129_ = _2034_ | _0598_;
  assign _0131_ = _2035_ | _0601_;
  assign _0133_ = _2036_ | _0604_;
  assign _0135_ = _2037_ | _0607_;
  assign _0137_ = _2038_ | _0610_;
  assign _0139_ = _2039_ | _0613_;
  assign _0141_ = _2040_ | _0616_;
  assign _0143_ = _2041_ | _0619_;
  assign _0145_ = _2042_ | _0622_;
  assign \gen_trigger_regs.tselect_we_t0  = _2043_ | _0625_;
  assign \gen_trigger_regs.tmatch_control_we_t0  = _2044_ | _0628_;
  assign _0147_ = _2045_ | _0631_;
  assign _0149_ = _2046_ | _0634_;
  assign \gen_trigger_regs.tmatch_value_we_t0  = _2047_ | _0637_;
  assign trigger_match_o_t0 = _2048_ | _0640_;
  assign _0517_ = | csr_addr_i_t0[11:10];
  assign _0518_ = | { \gen_trigger_regs.selected_tmatch_value_t0 , pc_if_i_t0 };
  assign _0521_ = | csr_op_i_t0;
  assign _0525_ = | csr_addr_i_t0[4:0];
  assign _0524_ = | csr_addr_i_t0;
  assign _2584_ = pc_if_i_t0 | \gen_trigger_regs.selected_tmatch_value_t0 ;
  assign _0336_ = ~ csr_addr_i_t0[11:10];
  assign _0337_ = ~ _2584_;
  assign _0344_ = ~ csr_wdata_int_t0[12:11];
  assign _0345_ = ~ csr_wdata_int_t0[1:0];
  assign _0359_ = ~ csr_op_i_t0;
  assign _0406_ = ~ csr_addr_i_t0[4:0];
  assign _0405_ = ~ csr_addr_i_t0;
  assign _1493_ = csr_addr_i[11:10] & _0336_;
  assign _1495_ = pc_if_i & _0337_;
  assign _1512_ = csr_wdata_int[12:11] & _0344_;
  assign _1514_ = csr_wdata_int[1:0] & _0345_;
  assign _1533_ = csr_op_i & _0359_;
  assign _1817_ = csr_addr_i[4:0] & _0406_;
  assign _1814_ = csr_addr_i & _0405_;
  assign _1494_ = 2'h3 & _0336_;
  assign _1496_ = \gen_trigger_regs.selected_tmatch_value  & _0337_;
  assign _1513_ = 2'h3 & _0344_;
  assign _1515_ = 2'h3 & _0345_;
  assign _1534_ = 2'h3 & _0359_;
  assign _1535_ = 2'h2 & _0359_;
  assign _1536_ = 2'h1 & _0359_;
  assign _1815_ = 12'h344 & _0405_;
  assign _1816_ = 12'h304 & _0405_;
  assign _1818_ = 5'h1f & _0406_;
  assign _1819_ = 5'h1e & _0406_;
  assign _1820_ = 5'h1d & _0406_;
  assign _1821_ = 5'h1c & _0406_;
  assign _1822_ = 5'h1b & _0406_;
  assign _1823_ = 5'h1a & _0406_;
  assign _1824_ = 5'h19 & _0406_;
  assign _1825_ = 5'h18 & _0406_;
  assign _1826_ = 5'h17 & _0406_;
  assign _1827_ = 5'h16 & _0406_;
  assign _1828_ = 5'h15 & _0406_;
  assign _1829_ = 5'h14 & _0406_;
  assign _1830_ = 5'h13 & _0406_;
  assign _1831_ = 5'h12 & _0406_;
  assign _1832_ = 5'h11 & _0406_;
  assign _1833_ = 5'h10 & _0406_;
  assign _1834_ = 5'h0f & _0406_;
  assign _1835_ = 5'h0e & _0406_;
  assign _1836_ = 5'h0d & _0406_;
  assign _1837_ = 5'h0c & _0406_;
  assign _1838_ = 5'h0b & _0406_;
  assign _1839_ = 5'h0a & _0406_;
  assign _1840_ = 5'h09 & _0406_;
  assign _1841_ = 5'h08 & _0406_;
  assign _1842_ = 5'h07 & _0406_;
  assign _1843_ = 5'h06 & _0406_;
  assign _1844_ = 5'h05 & _0406_;
  assign _1845_ = 5'h04 & _0406_;
  assign _1846_ = 5'h03 & _0406_;
  assign _1847_ = 5'h02 & _0406_;
  assign _1848_ = 5'h01 & _0406_;
  assign _1849_ = 12'h342 & _0405_;
  assign _1850_ = 12'h320 & _0405_;
  assign _1851_ = 12'h7b3 & _0405_;
  assign _1852_ = 12'h7b2 & _0405_;
  assign _1853_ = 12'h7b1 & _0405_;
  assign _1854_ = 12'h7b0 & _0405_;
  assign _1855_ = 12'h3bf & _0405_;
  assign _1856_ = 12'h3be & _0405_;
  assign _1857_ = 12'h3bd & _0405_;
  assign _1858_ = 12'h3bc & _0405_;
  assign _1859_ = 12'h3bb & _0405_;
  assign _1860_ = 12'h3ba & _0405_;
  assign _1861_ = 12'h3b9 & _0405_;
  assign _1862_ = 12'h3b8 & _0405_;
  assign _1863_ = 12'h3b7 & _0405_;
  assign _1864_ = 12'h3b6 & _0405_;
  assign _1865_ = 12'h3b5 & _0405_;
  assign _1866_ = 12'h3b4 & _0405_;
  assign _1867_ = 12'h3b3 & _0405_;
  assign _1868_ = 12'h3b2 & _0405_;
  assign _1869_ = 12'h3b1 & _0405_;
  assign _1870_ = 12'h3b0 & _0405_;
  assign _1871_ = 12'h3a3 & _0405_;
  assign _1872_ = 12'h3a2 & _0405_;
  assign _1873_ = 12'h3a1 & _0405_;
  assign _1874_ = 12'h3a0 & _0405_;
  assign _1875_ = 12'h343 & _0405_;
  assign _1876_ = 12'h341 & _0405_;
  assign _1877_ = 12'h305 & _0405_;
  assign _1878_ = 12'h340 & _0405_;
  assign _1879_ = 12'h301 & _0405_;
  assign _1880_ = 12'h300 & _0405_;
  assign _1881_ = 12'hf14 & _0405_;
  assign _1883_ = 12'hb13 & _0405_;
  assign _1884_ = 12'hb14 & _0405_;
  assign _1885_ = 12'hb15 & _0405_;
  assign _1886_ = 12'hb16 & _0405_;
  assign _1887_ = 12'hb17 & _0405_;
  assign _1888_ = 12'hb18 & _0405_;
  assign _1889_ = 12'hb19 & _0405_;
  assign _1890_ = 12'hb1a & _0405_;
  assign _1891_ = 12'hb1b & _0405_;
  assign _1892_ = 12'hb1c & _0405_;
  assign _1893_ = 12'hb1d & _0405_;
  assign _1894_ = 12'hb1e & _0405_;
  assign _1895_ = 12'hb1f & _0405_;
  assign _1896_ = 12'h323 & _0405_;
  assign _1897_ = 12'h324 & _0405_;
  assign _1898_ = 12'h32d & _0405_;
  assign _1899_ = 12'h32e & _0405_;
  assign _1900_ = 12'h32f & _0405_;
  assign _1901_ = 12'h330 & _0405_;
  assign _1902_ = 12'h331 & _0405_;
  assign _1903_ = 12'h332 & _0405_;
  assign _1904_ = 12'h333 & _0405_;
  assign _1905_ = 12'h334 & _0405_;
  assign _1906_ = 12'h335 & _0405_;
  assign _1907_ = 12'h336 & _0405_;
  assign _1908_ = 12'h325 & _0405_;
  assign _1909_ = 12'h337 & _0405_;
  assign _1910_ = 12'h338 & _0405_;
  assign _1911_ = 12'h339 & _0405_;
  assign _1912_ = 12'h33a & _0405_;
  assign _1913_ = 12'h33b & _0405_;
  assign _1914_ = 12'h33c & _0405_;
  assign _1915_ = 12'h33d & _0405_;
  assign _1916_ = 12'h33e & _0405_;
  assign _1917_ = 12'h33f & _0405_;
  assign _1918_ = 12'h326 & _0405_;
  assign _1919_ = 12'h327 & _0405_;
  assign _1920_ = 12'h328 & _0405_;
  assign _1921_ = 12'h329 & _0405_;
  assign _1922_ = 12'h32a & _0405_;
  assign _1923_ = 12'h32b & _0405_;
  assign _1924_ = 12'h32c & _0405_;
  assign _1925_ = 12'h7c1 & _0405_;
  assign _1926_ = 12'h7c0 & _0405_;
  assign _1927_ = 12'h7aa & _0405_;
  assign _1928_ = 12'h7a8 & _0405_;
  assign _1929_ = 12'h7a3 & _0405_;
  assign _1930_ = 12'h7a2 & _0405_;
  assign _1931_ = 12'h7a1 & _0405_;
  assign _1932_ = 12'h7a0 & _0405_;
  assign _1933_ = 12'hb80 & _0405_;
  assign _1934_ = 12'hb82 & _0405_;
  assign _1935_ = 12'hb8b & _0405_;
  assign _1936_ = 12'hb8c & _0405_;
  assign _1937_ = 12'hb8d & _0405_;
  assign _1938_ = 12'hb8e & _0405_;
  assign _1939_ = 12'hb8f & _0405_;
  assign _1940_ = 12'hb90 & _0405_;
  assign _1941_ = 12'hb91 & _0405_;
  assign _1942_ = 12'hb92 & _0405_;
  assign _1943_ = 12'hb93 & _0405_;
  assign _1944_ = 12'hb94 & _0405_;
  assign _1945_ = 12'hb83 & _0405_;
  assign _1946_ = 12'hb95 & _0405_;
  assign _1947_ = 12'hb96 & _0405_;
  assign _1948_ = 12'hb97 & _0405_;
  assign _1949_ = 12'hb98 & _0405_;
  assign _1950_ = 12'hb99 & _0405_;
  assign _1951_ = 12'hb9a & _0405_;
  assign _1952_ = 12'hb9b & _0405_;
  assign _1953_ = 12'hb9c & _0405_;
  assign _1954_ = 12'hb9d & _0405_;
  assign _1955_ = 12'hb9e & _0405_;
  assign _1956_ = 12'hb84 & _0405_;
  assign _1957_ = 12'hb9f & _0405_;
  assign _1958_ = 12'hb85 & _0405_;
  assign _1959_ = 12'hb86 & _0405_;
  assign _1960_ = 12'hb87 & _0405_;
  assign _1961_ = 12'hb88 & _0405_;
  assign _1962_ = 12'hb89 & _0405_;
  assign _1963_ = 12'hb8a & _0405_;
  assign _1964_ = 12'hb00 & _0405_;
  assign _1965_ = 12'hb02 & _0405_;
  assign _1966_ = 12'hb0b & _0405_;
  assign _1967_ = 12'hb0c & _0405_;
  assign _1968_ = 12'hb0d & _0405_;
  assign _1969_ = 12'hb0e & _0405_;
  assign _1970_ = 12'hb0f & _0405_;
  assign _1971_ = 12'hb10 & _0405_;
  assign _1972_ = 12'hb11 & _0405_;
  assign _1973_ = 12'hb12 & _0405_;
  assign _1974_ = 12'hb03 & _0405_;
  assign _1975_ = 12'hb04 & _0405_;
  assign _1976_ = 12'hb05 & _0405_;
  assign _1977_ = 12'hb06 & _0405_;
  assign _1978_ = 12'hb07 & _0405_;
  assign _1979_ = 12'hb08 & _0405_;
  assign _1980_ = 12'hb09 & _0405_;
  assign _1981_ = 12'hb0a & _0405_;
  assign _1982_ = 12'h306 & _0405_;
  assign _3068_ = _1493_ == _1494_;
  assign _3069_ = _1495_ == _1496_;
  assign _3070_ = _1512_ == _1513_;
  assign _3071_ = _1514_ == _1515_;
  assign _3072_ = _1533_ == _1534_;
  assign _3073_ = _1533_ == _1535_;
  assign _3074_ = _1533_ == _1536_;
  assign _3075_ = _1814_ == _1815_;
  assign _3076_ = _1814_ == _1816_;
  assign _3077_ = _1817_ == _1818_;
  assign _3078_ = _1817_ == _1819_;
  assign _3079_ = _1817_ == _1820_;
  assign _3080_ = _1817_ == _1821_;
  assign _3081_ = _1817_ == _1822_;
  assign _3082_ = _1817_ == _1823_;
  assign _3083_ = _1817_ == _1824_;
  assign _3084_ = _1817_ == _1825_;
  assign _3085_ = _1817_ == _1826_;
  assign _3086_ = _1817_ == _1827_;
  assign _3087_ = _1817_ == _1828_;
  assign _3088_ = _1817_ == _1829_;
  assign _3089_ = _1817_ == _1830_;
  assign _3090_ = _1817_ == _1831_;
  assign _3091_ = _1817_ == _1832_;
  assign _3092_ = _1817_ == _1833_;
  assign _3093_ = _1817_ == _1834_;
  assign _3094_ = _1817_ == _1835_;
  assign _3095_ = _1817_ == _1836_;
  assign _3096_ = _1817_ == _1837_;
  assign _3097_ = _1817_ == _1838_;
  assign _3098_ = _1817_ == _1839_;
  assign _3099_ = _1817_ == _1840_;
  assign _3100_ = _1817_ == _1841_;
  assign _3101_ = _1817_ == _1842_;
  assign _3102_ = _1817_ == _1843_;
  assign _3103_ = _1817_ == _1844_;
  assign _3104_ = _1817_ == _1845_;
  assign _3105_ = _1817_ == _1846_;
  assign _3106_ = _1817_ == _1847_;
  assign _3107_ = _1817_ == _1848_;
  assign _3108_ = _1814_ == _1849_;
  assign _3109_ = _1814_ == _1850_;
  assign _3110_ = _1814_ == _1851_;
  assign _3111_ = _1814_ == _1852_;
  assign _3112_ = _1814_ == _1853_;
  assign _3113_ = _1814_ == _1854_;
  assign _3114_ = _1814_ == _1855_;
  assign _3115_ = _1814_ == _1856_;
  assign _3116_ = _1814_ == _1857_;
  assign _3117_ = _1814_ == _1858_;
  assign _3118_ = _1814_ == _1859_;
  assign _3119_ = _1814_ == _1860_;
  assign _3120_ = _1814_ == _1861_;
  assign _3121_ = _1814_ == _1862_;
  assign _3122_ = _1814_ == _1863_;
  assign _3123_ = _1814_ == _1864_;
  assign _3124_ = _1814_ == _1865_;
  assign _3125_ = _1814_ == _1866_;
  assign _3126_ = _1814_ == _1867_;
  assign _3127_ = _1814_ == _1868_;
  assign _3128_ = _1814_ == _1869_;
  assign _3129_ = _1814_ == _1870_;
  assign _3130_ = _1814_ == _1871_;
  assign _3131_ = _1814_ == _1872_;
  assign _3132_ = _1814_ == _1873_;
  assign _3133_ = _1814_ == _1874_;
  assign _3134_ = _1814_ == _1875_;
  assign _3135_ = _1814_ == _1876_;
  assign _3136_ = _1814_ == _1877_;
  assign _3137_ = _1814_ == _1878_;
  assign _3138_ = _1814_ == _1879_;
  assign _3139_ = _1814_ == _1880_;
  assign _3140_ = _1814_ == _1881_;
  assign _3141_ = _1814_ == _1883_;
  assign _3142_ = _1814_ == _1884_;
  assign _3143_ = _1814_ == _1885_;
  assign _3144_ = _1814_ == _1886_;
  assign _3145_ = _1814_ == _1887_;
  assign _3146_ = _1814_ == _1888_;
  assign _3147_ = _1814_ == _1889_;
  assign _3148_ = _1814_ == _1890_;
  assign _3149_ = _1814_ == _1891_;
  assign _3150_ = _1814_ == _1892_;
  assign _3151_ = _1814_ == _1893_;
  assign _3152_ = _1814_ == _1894_;
  assign _3153_ = _1814_ == _1895_;
  assign _3154_ = _1814_ == _1896_;
  assign _3155_ = _1814_ == _1897_;
  assign _3156_ = _1814_ == _1898_;
  assign _3157_ = _1814_ == _1899_;
  assign _3158_ = _1814_ == _1900_;
  assign _3159_ = _1814_ == _1901_;
  assign _3160_ = _1814_ == _1902_;
  assign _3161_ = _1814_ == _1903_;
  assign _3162_ = _1814_ == _1904_;
  assign _3163_ = _1814_ == _1905_;
  assign _3164_ = _1814_ == _1906_;
  assign _3165_ = _1814_ == _1907_;
  assign _3166_ = _1814_ == _1908_;
  assign _3167_ = _1814_ == _1909_;
  assign _3168_ = _1814_ == _1910_;
  assign _3169_ = _1814_ == _1911_;
  assign _3170_ = _1814_ == _1912_;
  assign _3171_ = _1814_ == _1913_;
  assign _3172_ = _1814_ == _1914_;
  assign _3173_ = _1814_ == _1915_;
  assign _3174_ = _1814_ == _1916_;
  assign _3175_ = _1814_ == _1917_;
  assign _3176_ = _1814_ == _1918_;
  assign _3177_ = _1814_ == _1919_;
  assign _3178_ = _1814_ == _1920_;
  assign _3179_ = _1814_ == _1921_;
  assign _3180_ = _1814_ == _1922_;
  assign _3181_ = _1814_ == _1923_;
  assign _3182_ = _1814_ == _1924_;
  assign _3183_ = _1814_ == _1925_;
  assign _3184_ = _1814_ == _1926_;
  assign _3185_ = _1814_ == _1927_;
  assign _3186_ = _1814_ == _1928_;
  assign _3187_ = _1814_ == _1929_;
  assign _3188_ = _1814_ == _1930_;
  assign _3189_ = _1814_ == _1931_;
  assign _3190_ = _1814_ == _1932_;
  assign _3191_ = _1814_ == _1933_;
  assign _3192_ = _1814_ == _1934_;
  assign _3193_ = _1814_ == _1935_;
  assign _3194_ = _1814_ == _1936_;
  assign _3195_ = _1814_ == _1937_;
  assign _3196_ = _1814_ == _1938_;
  assign _3197_ = _1814_ == _1939_;
  assign _3198_ = _1814_ == _1940_;
  assign _3199_ = _1814_ == _1941_;
  assign _3200_ = _1814_ == _1942_;
  assign _3201_ = _1814_ == _1943_;
  assign _3202_ = _1814_ == _1944_;
  assign _3203_ = _1814_ == _1945_;
  assign _3204_ = _1814_ == _1946_;
  assign _3205_ = _1814_ == _1947_;
  assign _3206_ = _1814_ == _1948_;
  assign _3207_ = _1814_ == _1949_;
  assign _3208_ = _1814_ == _1950_;
  assign _3209_ = _1814_ == _1951_;
  assign _3210_ = _1814_ == _1952_;
  assign _3211_ = _1814_ == _1953_;
  assign _3212_ = _1814_ == _1954_;
  assign _3213_ = _1814_ == _1955_;
  assign _3214_ = _1814_ == _1956_;
  assign _3215_ = _1814_ == _1957_;
  assign _3216_ = _1814_ == _1958_;
  assign _3217_ = _1814_ == _1959_;
  assign _3218_ = _1814_ == _1960_;
  assign _3219_ = _1814_ == _1961_;
  assign _3220_ = _1814_ == _1962_;
  assign _3221_ = _1814_ == _1963_;
  assign _3222_ = _1814_ == _1964_;
  assign _3223_ = _1814_ == _1965_;
  assign _3224_ = _1814_ == _1966_;
  assign _3225_ = _1814_ == _1967_;
  assign _3226_ = _1814_ == _1968_;
  assign _3227_ = _1814_ == _1969_;
  assign _3228_ = _1814_ == _1970_;
  assign _3229_ = _1814_ == _1971_;
  assign _3230_ = _1814_ == _1972_;
  assign _3231_ = _1814_ == _1973_;
  assign _3232_ = _1814_ == _1974_;
  assign _3233_ = _1814_ == _1975_;
  assign _3234_ = _1814_ == _1976_;
  assign _3235_ = _1814_ == _1977_;
  assign _3236_ = _1814_ == _1978_;
  assign _3237_ = _1814_ == _1979_;
  assign _3238_ = _1814_ == _1980_;
  assign _3239_ = _1814_ == _1981_;
  assign _3240_ = _1814_ == _1982_;
  assign _3730_ = _3068_ & _0517_;
  assign _3745_ = _3069_ & _0518_;
  assign _3753_ = _3070_ & _0519_;
  assign _3757_ = _3071_ & _0520_;
  assign _3732_ = _3072_ & _0521_;
  assign _3734_ = _3073_ & _0521_;
  assign _3736_ = _3074_ & _0521_;
  assign _3893_ = _3075_ & _0524_;
  assign _0051_ = _3076_ & _0524_;
  assign _3895_ = _3077_ & _0525_;
  assign _3897_ = _3078_ & _0525_;
  assign _3899_ = _3079_ & _0525_;
  assign _3901_ = _3080_ & _0525_;
  assign _3903_ = _3081_ & _0525_;
  assign _3905_ = _3082_ & _0525_;
  assign _3907_ = _3083_ & _0525_;
  assign _3909_ = _3084_ & _0525_;
  assign _3911_ = _3085_ & _0525_;
  assign _3913_ = _3086_ & _0525_;
  assign _3915_ = _3087_ & _0525_;
  assign _3917_ = _3088_ & _0525_;
  assign _3919_ = _3089_ & _0525_;
  assign _3921_ = _3090_ & _0525_;
  assign _3923_ = _3091_ & _0525_;
  assign _3925_ = _3092_ & _0525_;
  assign _3927_ = _3093_ & _0525_;
  assign _3929_ = _3094_ & _0525_;
  assign _3931_ = _3095_ & _0525_;
  assign _3933_ = _3096_ & _0525_;
  assign _3935_ = _3097_ & _0525_;
  assign _3937_ = _3098_ & _0525_;
  assign _3939_ = _3099_ & _0525_;
  assign _3941_ = _3100_ & _0525_;
  assign _3943_ = _3101_ & _0525_;
  assign _3945_ = _3102_ & _0525_;
  assign _3947_ = _3103_ & _0525_;
  assign _3949_ = _3104_ & _0525_;
  assign _3951_ = _3105_ & _0525_;
  assign _3953_ = _3106_ & _0525_;
  assign _3955_ = _3107_ & _0525_;
  assign _0039_ = _3108_ & _0524_;
  assign _0041_ = _3109_ & _0524_;
  assign _0033_ = _3110_ & _0524_;
  assign _0031_ = _3111_ & _0524_;
  assign _0029_ = _3112_ & _0524_;
  assign _0025_ = _3113_ & _0524_;
  assign _3849_ = _3114_ & _0524_;
  assign _3851_ = _3115_ & _0524_;
  assign _3853_ = _3116_ & _0524_;
  assign _3855_ = _3117_ & _0524_;
  assign _3857_ = _3118_ & _0524_;
  assign _3859_ = _3119_ & _0524_;
  assign _3861_ = _3120_ & _0524_;
  assign _3863_ = _3121_ & _0524_;
  assign _3865_ = _3122_ & _0524_;
  assign _3867_ = _3123_ & _0524_;
  assign _3869_ = _3124_ & _0524_;
  assign _3871_ = _3125_ & _0524_;
  assign _3873_ = _3126_ & _0524_;
  assign _3875_ = _3127_ & _0524_;
  assign _3877_ = _3128_ & _0524_;
  assign _3879_ = _3129_ & _0524_;
  assign _3881_ = _3130_ & _0524_;
  assign _3883_ = _3131_ & _0524_;
  assign _3885_ = _3132_ & _0524_;
  assign _3887_ = _3133_ & _0524_;
  assign _0063_ = _3134_ & _0524_;
  assign _0045_ = _3135_ & _0524_;
  assign _3838_ = _3136_ & _0524_;
  assign _0053_ = _3137_ & _0524_;
  assign _3891_ = _3138_ & _0524_;
  assign _0059_ = _3139_ & _0524_;
  assign _3889_ = _3140_ & _0524_;
  assign _3829_[18] = _3141_ & _0524_;
  assign _3829_[19] = _3142_ & _0524_;
  assign _3829_[20] = _3143_ & _0524_;
  assign _3829_[21] = _3144_ & _0524_;
  assign _3829_[22] = _3145_ & _0524_;
  assign _3829_[23] = _3146_ & _0524_;
  assign _3829_[24] = _3147_ & _0524_;
  assign _3829_[25] = _3148_ & _0524_;
  assign _3829_[26] = _3149_ & _0524_;
  assign _3829_[27] = _3150_ & _0524_;
  assign _3829_[28] = _3151_ & _0524_;
  assign _3829_[29] = _3152_ & _0524_;
  assign _3829_[30] = _3153_ & _0524_;
  assign _3845_[0] = _3154_ & _0524_;
  assign _3845_[1] = _3155_ & _0524_;
  assign _3845_[10] = _3156_ & _0524_;
  assign _3845_[11] = _3157_ & _0524_;
  assign _3845_[12] = _3158_ & _0524_;
  assign _3845_[13] = _3159_ & _0524_;
  assign _3845_[14] = _3160_ & _0524_;
  assign _3845_[15] = _3161_ & _0524_;
  assign _3845_[16] = _3162_ & _0524_;
  assign _3845_[17] = _3163_ & _0524_;
  assign _3845_[18] = _3164_ & _0524_;
  assign _3845_[19] = _3165_ & _0524_;
  assign _3845_[2] = _3166_ & _0524_;
  assign _3845_[20] = _3167_ & _0524_;
  assign _3845_[21] = _3168_ & _0524_;
  assign _3845_[22] = _3169_ & _0524_;
  assign _3845_[23] = _3170_ & _0524_;
  assign _3845_[24] = _3171_ & _0524_;
  assign _3845_[25] = _3172_ & _0524_;
  assign _3845_[26] = _3173_ & _0524_;
  assign _3845_[27] = _3174_ & _0524_;
  assign _3845_[28] = _3175_ & _0524_;
  assign _3845_[3] = _3176_ & _0524_;
  assign _3845_[4] = _3177_ & _0524_;
  assign _3845_[5] = _3178_ & _0524_;
  assign _3845_[6] = _3179_ & _0524_;
  assign _3845_[7] = _3180_ & _0524_;
  assign _3845_[8] = _3181_ & _0524_;
  assign _3845_[9] = _3182_ & _0524_;
  assign _3957_ = _3183_ & _0524_;
  assign _0021_ = _3184_ & _0524_;
  assign _3959_ = _3185_ & _0524_;
  assign _3961_ = _3186_ & _0524_;
  assign _3963_ = _3187_ & _0524_;
  assign _3743_ = _3188_ & _0524_;
  assign _3741_ = _3189_ & _0524_;
  assign _3738_ = _3190_ & _0524_;
  assign _3825_[0] = _3191_ & _0524_;
  assign _3825_[1] = _3192_ & _0524_;
  assign _3825_[10] = _3193_ & _0524_;
  assign _3825_[11] = _3194_ & _0524_;
  assign _3825_[12] = _3195_ & _0524_;
  assign _3825_[13] = _3196_ & _0524_;
  assign _3825_[14] = _3197_ & _0524_;
  assign _3825_[15] = _3198_ & _0524_;
  assign _3825_[16] = _3199_ & _0524_;
  assign _3825_[17] = _3200_ & _0524_;
  assign _3825_[18] = _3201_ & _0524_;
  assign _3825_[19] = _3202_ & _0524_;
  assign _3825_[2] = _3203_ & _0524_;
  assign _3825_[20] = _3204_ & _0524_;
  assign _3825_[21] = _3205_ & _0524_;
  assign _3825_[22] = _3206_ & _0524_;
  assign _3825_[23] = _3207_ & _0524_;
  assign _3825_[24] = _3208_ & _0524_;
  assign _3825_[25] = _3209_ & _0524_;
  assign _3825_[26] = _3210_ & _0524_;
  assign _3825_[27] = _3211_ & _0524_;
  assign _3825_[28] = _3212_ & _0524_;
  assign _3825_[29] = _3213_ & _0524_;
  assign _3825_[3] = _3214_ & _0524_;
  assign _3825_[30] = _3215_ & _0524_;
  assign _3825_[4] = _3216_ & _0524_;
  assign _3825_[5] = _3217_ & _0524_;
  assign _3825_[6] = _3218_ & _0524_;
  assign _3825_[7] = _3219_ & _0524_;
  assign _3825_[8] = _3220_ & _0524_;
  assign _3825_[9] = _3221_ & _0524_;
  assign _3829_[0] = _3222_ & _0524_;
  assign _3829_[1] = _3223_ & _0524_;
  assign _3829_[10] = _3224_ & _0524_;
  assign _3829_[11] = _3225_ & _0524_;
  assign _3829_[12] = _3226_ & _0524_;
  assign _3829_[13] = _3227_ & _0524_;
  assign _3829_[14] = _3228_ & _0524_;
  assign _3829_[15] = _3229_ & _0524_;
  assign _3829_[16] = _3230_ & _0524_;
  assign _3829_[17] = _3231_ & _0524_;
  assign _3829_[2] = _3232_ & _0524_;
  assign _3829_[3] = _3233_ & _0524_;
  assign _3829_[4] = _3234_ & _0524_;
  assign _3829_[5] = _3235_ & _0524_;
  assign _3829_[6] = _3236_ & _0524_;
  assign _3829_[7] = _3237_ & _0524_;
  assign _3829_[8] = _3238_ & _0524_;
  assign _3829_[9] = _3239_ & _0524_;
  assign _3965_ = _3240_ & _0524_;
  reg [11:0] _4657_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) _4657_ <= 12'h000;
    else if (mcountinhibit_we) _4657_ <= { csr_wdata_int[12:2], csr_wdata_int[0] };
  assign { mcountinhibit[12:2], mcountinhibit[0] } = _4657_;
  assign _0150_ = { _1497_, _1499_ } > { _2586_, _2588_ };
  assign _0151_ = { _2585_, _2587_ } > { _1498_, _1500_ };
  assign illegal_csr_priv_t0 = _0150_ ^ _0151_;
  assign _0338_ = ~ csr_addr_i_t0[8];
  assign _0339_ = ~ csr_addr_i_t0[9];
  assign _0340_ = ~ priv_mode_id_o_t0[0];
  assign _0341_ = ~ priv_mode_id_o_t0[1];
  assign _1497_ = csr_addr_i[9] & _0339_;
  assign _1498_ = priv_mode_id_o[1] & _0341_;
  assign _2585_ = csr_addr_i[9] | csr_addr_i_t0[9];
  assign _2586_ = priv_mode_id_o[1] | priv_mode_id_o_t0[1];
  assign _1499_ = csr_addr_i[8] & _0338_;
  assign _1500_ = priv_mode_id_o[0] & _0340_;
  assign _2587_ = csr_addr_i[8] | csr_addr_i_t0[8];
  assign _2588_ = priv_mode_id_o[0] | priv_mode_id_o_t0[0];
  assign _1501_ = _3730_ & csr_wr;
  assign _1504_ = _3753_ & _3754_;
  assign _1507_ = _3757_ & _3758_;
  assign _1502_ = csr_wr_t0 & _3729_;
  assign _1505_ = _3755_ & _3752_;
  assign _1508_ = _3759_ & _3756_;
  assign _1503_ = _3730_ & csr_wr_t0;
  assign _1506_ = _3753_ & _3755_;
  assign _1509_ = _3757_ & _3759_;
  assign _2589_ = _1501_ | _1502_;
  assign _2590_ = _1504_ | _1505_;
  assign _2591_ = _1507_ | _1508_;
  assign illegal_csr_write_t0 = _2589_ | _1503_;
  assign _3747_ = _2590_ | _1506_;
  assign _3749_ = _2591_ | _1509_;
  assign _0484_ = | { _0051_, _0053_, _0045_, _0039_, _0063_, _0041_, _0021_, _0059_, _3965_, _3963_, _3961_, _3959_, _3957_, _3893_, _3891_, _3889_, _3887_, _3885_, _3883_, _3881_, _3879_, _3877_, _3875_, _3873_, _3871_, _3869_, _3867_, _3865_, _3863_, _3861_, _3859_, _3857_, _3855_, _3853_, _3851_, _3849_, _3845_, _3838_, _3829_, _3825_, _3743_, _3741_, _3738_ };
  assign _0485_ = | { _0025_, _0029_, _0031_, _0033_ };
  assign _0486_ = | { _3955_, _3931_, _3929_, _3927_, _3925_, _3923_, _3921_, _3919_, _3917_, _3915_, _3913_, _3911_, _3909_, _3907_, _3905_, _3903_, _3901_, _3899_, _3897_, _3895_ };
  assign _0487_ = | { _3736_, _3785_ };
  assign _0488_ = | { _3891_, _3741_ };
  assign _0489_ = | { _0045_, _0039_, _1998_ };
  assign _0490_ = | { _0045_, _1998_, _3838_ };
  assign _0491_ = | { _2008_, _3825_, _3741_ };
  assign _0492_ = | { _0039_, _0063_, _2012_ };
  assign _0493_ = | { _0031_, _0033_, _0041_, _2010_, _2008_, _3825_, _3741_ };
  assign _0494_ = | { _2008_, _3829_, _3825_, _3741_ };
  assign _0495_ = | { _0051_, _0053_, _3838_ };
  assign _0496_ = | { _0045_, _0039_, _0063_, _2020_ };
  assign _0497_ = | { _0029_, _0031_, _0033_, _2018_, _2008_, _3829_, _3825_, _3741_ };
  assign _0498_ = | { _3935_, _3933_, _3955_, _3931_, _3929_, _3927_, _3925_, _3923_, _3921_, _3919_, _3917_, _3915_, _3913_, _3911_, _3909_, _3907_, _3905_, _3903_, _3901_, _3899_, _3897_, _3895_ };
  assign _0499_ = | { _3947_, _3945_, _3943_ };
  assign _0500_ = | { _3941_, _3939_, _3937_, _3935_, _3933_, _3955_, _3931_, _3929_, _3927_, _3925_, _3923_, _3921_, _3919_, _3917_, _3915_, _3913_, _3911_, _3909_, _3907_, _3905_, _3903_, _3901_, _3899_, _3897_, _3895_ };
  assign _0501_ = | { _2022_, _3829_, _3825_ };
  assign _0502_ = | { _0045_, _0063_, _2020_, _3838_ };
  assign _0503_ = | { _0029_, _0031_, _0033_, _2018_, _2022_, _3829_, _3825_ };
  assign _0504_ = | { _3829_, _3825_, _3743_ };
  assign _0505_ = | { _0031_, _0033_, _2018_, _3829_, _3825_, _3743_ };
  assign _0506_ = | { _0025_, _0029_, _0031_, _1996_, _1994_, _3845_, _3829_ };
  assign _0507_ = | { _0045_, _0063_, _2020_ };
  assign _0508_ = | { _0029_, _0031_, _1996_, _1994_, _3845_, _3829_ };
  assign _0509_ = | { _1994_, _3845_, _3829_ };
  assign _0510_ = | { _0045_, _2004_, _3838_ };
  assign _0511_ = | { _2008_, _3825_, _3741_, _3738_ };
  assign _0512_ = | { _0045_, _0039_, _0063_, _2012_ };
  assign _0513_ = | { _0031_, _0033_, _0041_, _2010_, _2008_, _3825_, _3741_, _3738_ };
  assign _0514_ = | { _2024_, _3829_, _3825_ };
  assign _0515_ = | { _0045_, _0063_, _2012_ };
  assign _0516_ = | { _0031_, _0033_, _2018_, _2024_, _3829_, _3825_ };
  assign _0519_ = | csr_wdata_int_t0[12:11];
  assign _0520_ = | csr_wdata_int_t0[1:0];
  assign _0522_ = | _3825_;
  assign _0523_ = | _3845_;
  assign _0526_ = | _3829_;
  assign _0527_ = | { _3734_, _3732_, _3736_ };
  assign _0528_ = | irqs_o_t0;
  assign _0165_ = ~ { _3965_, _3963_, _3961_, _3959_, _3957_, _3893_, _3891_, _3889_, _3887_, _3885_, _3883_, _3881_, _3879_, _3877_, _3875_, _3873_, _3871_, _3869_, _3867_, _3865_, _3863_, _3861_, _3859_, _3857_, _3855_, _3853_, _3851_, _3849_, _3845_, _0051_, _0053_, _0045_, _0039_, _0063_, _3838_, _0041_, _0021_, _3829_, _3825_, _0059_, _3743_, _3741_, _3738_ };
  assign _0166_ = ~ { _0029_, _0031_, _0033_, _0025_ };
  assign _0167_ = ~ { _3955_, _3931_, _3929_, _3927_, _3925_, _3923_, _3921_, _3919_, _3917_, _3915_, _3913_, _3911_, _3909_, _3907_, _3905_, _3903_, _3901_, _3899_, _3897_, _3895_ };
  assign _0168_ = ~ { _3736_, _3785_ };
  assign _0169_ = ~ { _3891_, _3741_ };
  assign _0190_ = ~ { _1998_, _0045_, _0039_ };
  assign _0191_ = ~ { _1998_, _0045_, _3838_ };
  assign _0192_ = ~ { _3825_, _2008_, _3741_ };
  assign _0193_ = ~ { _0039_, _0063_, _2012_ };
  assign _0194_ = ~ { _0031_, _0033_, _0041_, _3825_, _2008_, _2010_, _3741_ };
  assign _0195_ = ~ { _3829_, _3825_, _2008_, _3741_ };
  assign _0196_ = ~ { _0051_, _0053_, _3838_ };
  assign _0197_ = ~ { _0045_, _0039_, _0063_, _2020_ };
  assign _0198_ = ~ { _0029_, _0031_, _0033_, _3829_, _3825_, _2008_, _3741_, _2018_ };
  assign _0199_ = ~ { _3955_, _3935_, _3933_, _3931_, _3929_, _3927_, _3925_, _3923_, _3921_, _3919_, _3917_, _3915_, _3913_, _3911_, _3909_, _3907_, _3905_, _3903_, _3901_, _3899_, _3897_, _3895_ };
  assign _0200_ = ~ { _3947_, _3945_, _3943_ };
  assign _0201_ = ~ { _3955_, _3941_, _3939_, _3937_, _3935_, _3933_, _3931_, _3929_, _3927_, _3925_, _3923_, _3921_, _3919_, _3917_, _3915_, _3913_, _3911_, _3909_, _3907_, _3905_, _3903_, _3901_, _3899_, _3897_, _3895_ };
  assign _0202_ = ~ { _2022_, _3829_, _3825_ };
  assign _0203_ = ~ { _0045_, _0063_, _3838_, _2020_ };
  assign _0204_ = ~ { _2022_, _0029_, _0031_, _0033_, _3829_, _3825_, _2018_ };
  assign _0205_ = ~ { _3829_, _3825_, _3743_ };
  assign _0206_ = ~ { _0031_, _0033_, _3829_, _3825_, _3743_, _2018_ };
  assign _0207_ = ~ { _1996_, _1994_, _3845_, _0029_, _0031_, _3829_, _0025_ };
  assign _0208_ = ~ { _0045_, _0063_, _2020_ };
  assign _0209_ = ~ { _1996_, _1994_, _3845_, _0029_, _0031_, _3829_ };
  assign _0210_ = ~ { _1994_, _3845_, _3829_ };
  assign _0211_ = ~ { _2004_, _0045_, _3838_ };
  assign _0212_ = ~ { _3825_, _2008_, _3741_, _3738_ };
  assign _0213_ = ~ { _0045_, _0039_, _0063_, _2012_ };
  assign _0214_ = ~ { _0031_, _0033_, _0041_, _3825_, _2008_, _2010_, _3741_, _3738_ };
  assign _0215_ = ~ { _3829_, _3825_, _2024_ };
  assign _0216_ = ~ { _0045_, _0063_, _2012_ };
  assign _0217_ = ~ { _0031_, _0033_, _3829_, _3825_, _2018_, _2024_ };
  assign _0403_ = ~ _3825_;
  assign _0404_ = ~ _3845_;
  assign _0407_ = ~ _3829_;
  assign _0408_ = ~ { _3736_, _3734_, _3732_ };
  assign _0409_ = ~ irqs_o_t0;
  assign _0644_ = { _3964_, _3962_, _3960_, _3958_, _3956_, _3892_, _3890_, _3888_, _3886_, _3884_, _3882_, _3880_, _3878_, _3876_, _3874_, _3872_, _3870_, _3868_, _3866_, _3864_, _3862_, _3860_, _3858_, _3856_, _3854_, _3852_, _3850_, _3848_, _3844_, _3843_, _3842_, _3841_, _3840_, _3839_, _3837_, _3833_, _3832_, _3828_, _3824_, _3823_, _3742_, _3740_, _3737_ } & _0165_;
  assign _0645_ = { _3836_, _3835_, _3834_, _3822_ } & _0166_;
  assign _0646_ = { _3954_, _3930_, _3928_, _3926_, _3924_, _3922_, _3920_, _3918_, _3916_, _3914_, _3912_, _3910_, _3908_, _3906_, _3904_, _3902_, _3900_, _3898_, _3896_, _3894_ } & _0167_;
  assign _0647_ = { _3735_, _3784_ } & _0168_;
  assign _0648_ = { _3890_, _3740_ } & _0169_;
  assign _0697_ = { _1997_, _3841_, _3840_ } & _0190_;
  assign _0698_ = { _1997_, _3841_, _3837_ } & _0191_;
  assign _0699_ = { _3824_, _2007_, _3740_ } & _0192_;
  assign _0700_ = { _3840_, _3839_, _2011_ } & _0193_;
  assign _0701_ = { _3835_, _3834_, _3833_, _3824_, _2007_, _2009_, _3740_ } & _0194_;
  assign _0702_ = { _3828_, _3824_, _2007_, _3740_ } & _0195_;
  assign _0703_ = { _3843_, _3842_, _3837_ } & _0196_;
  assign _0704_ = { _3841_, _3840_, _3839_, _2019_ } & _0197_;
  assign _0705_ = { _3836_, _3835_, _3834_, _3828_, _3824_, _2007_, _3740_, _2017_ } & _0198_;
  assign _0706_ = { _3954_, _3934_, _3932_, _3930_, _3928_, _3926_, _3924_, _3922_, _3920_, _3918_, _3916_, _3914_, _3912_, _3910_, _3908_, _3906_, _3904_, _3902_, _3900_, _3898_, _3896_, _3894_ } & _0199_;
  assign _0707_ = { _3946_, _3944_, _3942_ } & _0200_;
  assign _0708_ = { _3954_, _3940_, _3938_, _3936_, _3934_, _3932_, _3930_, _3928_, _3926_, _3924_, _3922_, _3920_, _3918_, _3916_, _3914_, _3912_, _3910_, _3908_, _3906_, _3904_, _3902_, _3900_, _3898_, _3896_, _3894_ } & _0201_;
  assign _0709_ = { _2021_, _3828_, _3824_ } & _0202_;
  assign _0710_ = { _3841_, _3839_, _3837_, _2019_ } & _0203_;
  assign _0711_ = { _2021_, _3836_, _3835_, _3834_, _3828_, _3824_, _2017_ } & _0204_;
  assign _0712_ = { _3828_, _3824_, _3742_ } & _0205_;
  assign _0713_ = { _3835_, _3834_, _3828_, _3824_, _3742_, _2017_ } & _0206_;
  assign _0714_ = { _1995_, _1993_, _3844_, _3836_, _3835_, _3828_, _3822_ } & _0207_;
  assign _0715_ = { _3841_, _3839_, _2019_ } & _0208_;
  assign _0716_ = { _1995_, _1993_, _3844_, _3836_, _3835_, _3828_ } & _0209_;
  assign _0717_ = { _1993_, _3844_, _3828_ } & _0210_;
  assign _0718_ = { _2003_, _3841_, _3837_ } & _0211_;
  assign _0719_ = { _3824_, _2007_, _3740_, _3737_ } & _0212_;
  assign _0720_ = { _3841_, _3840_, _3839_, _2011_ } & _0213_;
  assign _0721_ = { _3835_, _3834_, _3833_, _3824_, _2007_, _2009_, _3740_, _3737_ } & _0214_;
  assign _0722_ = { _3828_, _3824_, _2023_ } & _0215_;
  assign _0723_ = { _3841_, _3839_, _2011_ } & _0216_;
  assign _0724_ = { _3835_, _3834_, _3828_, _3824_, _2017_, _2023_ } & _0217_;
  assign _1812_ = _3824_ & _0403_;
  assign _1813_ = _3844_ & _0404_;
  assign _1882_ = _3828_ & _0407_;
  assign _1983_ = { _3735_, _3733_, _3731_ } & _0408_;
  assign _1984_ = irqs_o & _0409_;
  assign _0530_ = ! _0644_;
  assign _0531_ = ! _0645_;
  assign _0532_ = ! _0646_;
  assign _0533_ = ! _0647_;
  assign _0534_ = ! _0648_;
  assign _0535_ = ! _0697_;
  assign _0536_ = ! _0698_;
  assign _0537_ = ! _0699_;
  assign _0538_ = ! _0700_;
  assign _0539_ = ! _0701_;
  assign _0540_ = ! _0702_;
  assign _0541_ = ! _0703_;
  assign _0542_ = ! _0704_;
  assign _0543_ = ! _0705_;
  assign _0544_ = ! _0706_;
  assign _0545_ = ! _0707_;
  assign _0546_ = ! _0708_;
  assign _0547_ = ! _0709_;
  assign _0548_ = ! _0710_;
  assign _0549_ = ! _0711_;
  assign _0550_ = ! _0712_;
  assign _0551_ = ! _0713_;
  assign _0552_ = ! _0714_;
  assign _0553_ = ! _0715_;
  assign _0554_ = ! _0716_;
  assign _0555_ = ! _0717_;
  assign _0556_ = ! _0718_;
  assign _0557_ = ! _0719_;
  assign _0558_ = ! _0720_;
  assign _0559_ = ! _0721_;
  assign _0560_ = ! _0722_;
  assign _0561_ = ! _0723_;
  assign _0562_ = ! _0724_;
  assign _0563_ = ! _1512_;
  assign _0564_ = ! _1514_;
  assign _0565_ = ! _1533_;
  assign _0566_ = ! _1812_;
  assign _0567_ = ! _1813_;
  assign _0568_ = ! _1882_;
  assign _0569_ = ! _1983_;
  assign _0570_ = ! _1984_;
  assign _0157_ = _0530_ & _0484_;
  assign _0159_ = _0531_ & _0485_;
  assign _0155_ = _0532_ & _0486_;
  assign _0161_ = _0533_ & _0487_;
  assign _0163_ = _0534_ & _0488_;
  assign _0431_ = _0535_ & _0489_;
  assign _0435_ = _0536_ & _0490_;
  assign _0441_ = _0537_ & _0491_;
  assign _0443_ = _0538_ & _0492_;
  assign _0445_ = _0539_ & _0493_;
  assign _0453_ = _0540_ & _0494_;
  assign _0455_ = _0541_ & _0495_;
  assign _0457_ = _0542_ & _0496_;
  assign _0459_ = _0543_ & _0497_;
  assign _0447_ = _0544_ & _0498_;
  assign _0449_ = _0545_ & _0499_;
  assign _0451_ = _0546_ & _0500_;
  assign _0461_ = _0547_ & _0501_;
  assign _0463_ = _0548_ & _0502_;
  assign _0465_ = _0549_ & _0503_;
  assign _0467_ = _0550_ & _0504_;
  assign _0471_ = _0551_ & _0505_;
  assign _0439_ = _0552_ & _0506_;
  assign _0473_ = _0553_ & _0507_;
  assign _0433_ = _0554_ & _0508_;
  assign _0429_ = _0555_ & _0509_;
  assign _0437_ = _0556_ & _0510_;
  assign _0475_ = _0557_ & _0511_;
  assign _0477_ = _0558_ & _0512_;
  assign _0479_ = _0559_ & _0513_;
  assign _0481_ = _0560_ & _0514_;
  assign _0469_ = _0561_ & _0515_;
  assign _0483_ = _0562_ & _0516_;
  assign _3755_ = _0563_ & _0519_;
  assign _3759_ = _0564_ & _0520_;
  assign _3785_ = _0565_ & _0521_;
  assign _3827_ = _0566_ & _0522_;
  assign _3847_ = _0567_ & _0523_;
  assign _3831_ = _0568_ & _0526_;
  assign csr_wr_t0 = _0569_ & _0527_;
  assign irq_pending_o_t0 = _0570_ & _0528_;
  assign _0152_ = { _1510_, _1511_ } < 32'd1;
  assign _0153_ = { _2592_, _2593_ } < 32'd1;
  assign _3751_ = _0152_ ^ _0153_;
  assign _0342_ = ~ csr_wdata_int_t0[30:0];
  assign _0343_ = ~ csr_wdata_int_t0[31];
  assign _1510_ = csr_wdata_int[31] & _0343_;
  assign _2592_ = csr_wdata_int[31] | csr_wdata_int_t0[31];
  assign _1511_ = csr_wdata_int[30:0] & _0342_;
  assign _2593_ = csr_wdata_int[30:0] | csr_wdata_int_t0[30:0];
  assign _0218_ = ~ { _3731_, _3731_, _3731_, _3731_, _3731_, _3731_, _3731_, _3731_, _3731_, _3731_, _3731_, _3731_, _3731_, _3731_, _3731_, _3731_, _3731_, _3731_, _3731_, _3731_, _3731_, _3731_, _3731_, _3731_, _3731_, _3731_, _3731_, _3731_, _3731_, _3731_, _3731_, _3731_ };
  assign _0219_ = ~ { _0160_, _0160_, _0160_, _0160_, _0160_, _0160_, _0160_, _0160_, _0160_, _0160_, _0160_, _0160_, _0160_, _0160_, _0160_, _0160_, _0160_, _0160_, _0160_, _0160_, _0160_, _0160_, _0160_, _0160_, _0160_, _0160_, _0160_, _0160_, _0160_, _0160_, _0160_, _0160_ };
  assign _0225_ = ~ _1997_;
  assign _0227_ = ~ _0430_;
  assign _0236_ = ~ { _3822_, _3822_, _3822_ };
  assign _0238_ = ~ { _1997_, _1997_, _1997_ };
  assign _0241_ = ~ { _2001_, _2001_, _2001_ };
  assign _0242_ = ~ { _0434_, _0434_, _0434_ };
  assign _0243_ = ~ { _0432_, _0432_, _0432_ };
  assign _0254_ = ~ { _0440_, _0440_, _0440_ };
  assign _0258_ = ~ { _2013_, _2013_, _2013_ };
  assign _0259_ = ~ { _0442_, _0442_, _0442_ };
  assign _0260_ = ~ { _0444_, _0444_, _0444_ };
  assign _0261_ = ~ { _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_ };
  assign _0262_ = ~ { _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_ };
  assign _0263_ = ~ { _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_ };
  assign _0264_ = ~ { _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_ };
  assign _0265_ = ~ { _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_ };
  assign _0266_ = ~ { _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_ };
  assign _0267_ = ~ { _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_ };
  assign _0268_ = ~ { _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_ };
  assign _0269_ = ~ { _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_ };
  assign _0270_ = ~ { _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_ };
  assign _0271_ = ~ { _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_ };
  assign _0272_ = ~ { _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_ };
  assign _0178_ = ~ _3740_;
  assign _0273_ = ~ _2007_;
  assign _0275_ = ~ _0452_;
  assign _0277_ = ~ _0454_;
  assign _0278_ = ~ _0456_;
  assign _0279_ = ~ _0458_;
  assign _0280_ = ~ { _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_ };
  assign _0281_ = ~ { _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_ };
  assign _0282_ = ~ { _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_ };
  assign _0283_ = ~ { _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_ };
  assign _0284_ = ~ { _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_ };
  assign _0285_ = ~ { _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_ };
  assign _0286_ = ~ { _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_ };
  assign _0287_ = ~ { _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_ };
  assign _0288_ = ~ { _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_ };
  assign _0289_ = ~ { _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_ };
  assign _0290_ = ~ { _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_ };
  assign _0291_ = ~ { _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_ };
  assign _0292_ = ~ { _3742_, _3742_, _3742_, _3742_, _3742_, _3742_, _3742_, _3742_, _3742_ };
  assign _0293_ = ~ { _3826_, _3826_, _3826_, _3826_, _3826_, _3826_, _3826_, _3826_, _3826_ };
  assign _0294_ = ~ { _2021_, _2021_, _2021_, _2021_, _2021_, _2021_, _2021_, _2021_, _2021_ };
  assign _0295_ = ~ { _3846_, _3846_, _3846_, _3846_, _3846_, _3846_, _3846_, _3846_, _3846_ };
  assign _0296_ = ~ { _3835_, _3835_, _3835_, _3835_, _3835_, _3835_, _3835_, _3835_, _3835_ };
  assign _0297_ = ~ { _3834_, _3834_, _3834_, _3834_, _3834_, _3834_, _3834_, _3834_, _3834_ };
  assign _0298_ = ~ { _2017_, _2017_, _2017_, _2017_, _2017_, _2017_, _2017_, _2017_, _2017_ };
  assign _0299_ = ~ { _0460_, _0460_, _0460_, _0460_, _0460_, _0460_, _0460_, _0460_, _0460_ };
  assign _0300_ = ~ { _3822_, _3822_, _3822_, _3822_, _3822_, _3822_, _3822_, _3822_, _3822_ };
  assign _0301_ = ~ { _3841_, _3841_, _3841_, _3841_, _3841_, _3841_, _3841_, _3841_, _3841_ };
  assign _0302_ = ~ { _3839_, _3839_, _3839_, _3839_, _3839_, _3839_, _3839_, _3839_, _3839_ };
  assign _0303_ = ~ { _2019_, _2019_, _2019_, _2019_, _2019_, _2019_, _2019_, _2019_, _2019_ };
  assign _0304_ = ~ { _3842_, _3842_, _3842_, _3842_, _3842_, _3842_, _3842_, _3842_, _3842_ };
  assign _0305_ = ~ { _3888_, _3888_, _3888_, _3888_, _3888_, _3888_, _3888_, _3888_, _3888_ };
  assign _0306_ = ~ { _3890_, _3890_, _3890_, _3890_, _3890_, _3890_, _3890_, _3890_, _3890_ };
  assign _0307_ = ~ { _2005_, _2005_, _2005_, _2005_, _2005_, _2005_, _2005_, _2005_, _2005_ };
  assign _0308_ = ~ { _0462_, _0462_, _0462_, _0462_, _0462_, _0462_, _0462_, _0462_, _0462_ };
  assign _0309_ = ~ { _0464_, _0464_, _0464_, _0464_, _0464_, _0464_, _0464_, _0464_, _0464_ };
  assign _0310_ = ~ { _3826_, _3826_, _3826_ };
  assign _0311_ = ~ { _3846_, _3846_, _3846_ };
  assign _0312_ = ~ { _2017_, _2017_, _2017_ };
  assign _0313_ = ~ { _0466_, _0466_, _0466_ };
  assign _0316_ = ~ { _0468_, _0468_, _0468_ };
  assign _0317_ = ~ { _0470_, _0470_, _0470_ };
  assign _0229_ = ~ { _3742_, _3742_, _3742_ };
  assign _0231_ = ~ { _1993_, _1993_, _1993_ };
  assign _0233_ = ~ { _3835_, _3835_, _3835_ };
  assign _0234_ = ~ { _1995_, _1995_, _1995_ };
  assign _0235_ = ~ { _0428_, _0428_, _0428_ };
  assign _0318_ = ~ { _3892_, _3892_, _3892_ };
  assign _0237_ = ~ { _3841_, _3841_, _3841_ };
  assign _0319_ = ~ { _2003_, _2003_, _2003_ };
  assign _0239_ = ~ { _3842_, _3842_, _3842_ };
  assign _0321_ = ~ { _2005_, _2005_, _2005_ };
  assign _0322_ = ~ { _0436_, _0436_, _0436_ };
  assign _0323_ = ~ { _0438_, _0438_, _0438_ };
  assign _0276_ = ~ _2019_;
  assign _0324_ = ~ _0472_;
  assign _0228_ = ~ _0432_;
  assign _0187_ = ~ _3830_;
  assign _0220_ = ~ _1993_;
  assign _0222_ = ~ _1995_;
  assign _0223_ = ~ _0428_;
  assign _0180_ = ~ _3892_;
  assign _0244_ = ~ _2003_;
  assign _0246_ = ~ _2005_;
  assign _0247_ = ~ _0436_;
  assign _0248_ = ~ _0438_;
  assign _0249_ = ~ { _3832_, _3832_, _3832_ };
  assign _0325_ = ~ { _3737_, _3737_, _3737_ };
  assign _0250_ = ~ { _3740_, _3740_, _3740_ };
  assign _0251_ = ~ { _2007_, _2007_, _2007_ };
  assign _0230_ = ~ { _3830_, _3830_, _3830_ };
  assign _0252_ = ~ { _3834_, _3834_, _3834_ };
  assign _0232_ = ~ { _3833_, _3833_, _3833_ };
  assign _0253_ = ~ { _2009_, _2009_, _2009_ };
  assign _0326_ = ~ { _0474_, _0474_, _0474_ };
  assign _0255_ = ~ { _3836_, _3836_, _3836_ };
  assign _0327_ = ~ { _3840_, _3840_, _3840_ };
  assign _0256_ = ~ { _3839_, _3839_, _3839_ };
  assign _0257_ = ~ { _2011_, _2011_, _2011_ };
  assign _0314_ = ~ { _3837_, _3837_, _3837_ };
  assign _0240_ = ~ { _3888_, _3888_, _3888_ };
  assign _0320_ = ~ { _3890_, _3890_, _3890_ };
  assign _0315_ = ~ { _1999_, _1999_, _1999_ };
  assign _0328_ = ~ { _0476_, _0476_, _0476_ };
  assign _0329_ = ~ { _0478_, _0478_, _0478_ };
  assign _0179_ = ~ _3742_;
  assign _0181_ = ~ _3826_;
  assign _0330_ = ~ _2023_;
  assign _0186_ = ~ _3846_;
  assign _0274_ = ~ _2017_;
  assign _0331_ = ~ _0480_;
  assign _0332_ = ~ _2011_;
  assign _0226_ = ~ _1999_;
  assign _0333_ = ~ _0468_;
  assign _0334_ = ~ _0482_;
  assign _0335_ = ~ _0156_;
  assign _0364_ = ~ { nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i };
  assign _0365_ = ~ { nmi_mode_i, nmi_mode_i };
  assign _0363_ = ~ nmi_mode_i;
  assign _0366_ = ~ { csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i };
  assign _0367_ = ~ { csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i };
  assign _0369_ = ~ { nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i };
  assign _0370_ = ~ { debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i };
  assign _0373_ = ~ { debug_mode_i, debug_mode_i };
  assign _0372_ = ~ { debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i };
  assign _0376_ = ~ { debug_csr_save_i, debug_csr_save_i, debug_csr_save_i };
  assign _0377_ = ~ { debug_csr_save_i, debug_csr_save_i };
  assign _0378_ = ~ { debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i };
  assign _0375_ = ~ { debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i };
  assign _0374_ = ~ debug_csr_save_i;
  assign _0379_ = ~ { debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i };
  assign _0380_ = ~ { csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i };
  assign _0381_ = ~ { csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i };
  assign _0382_ = ~ { csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i };
  assign _0368_ = ~ { csr_save_cause_i, csr_save_cause_i, csr_save_cause_i };
  assign _0385_ = ~ { csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i };
  assign _0386_ = ~ { csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i };
  assign _0387_ = ~ { csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i };
  assign _0388_ = ~ { csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i };
  assign _0389_ = ~ { csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i };
  assign _0383_ = ~ { csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i };
  assign _0360_ = ~ csr_restore_mret_i;
  assign _0361_ = ~ csr_restore_dret_i;
  assign _0362_ = ~ csr_save_cause_i;
  assign _0371_ = ~ debug_mode_i;
  assign _0390_ = ~ { csr_restore_mret_i, csr_restore_mret_i };
  assign _0391_ = ~ { csr_restore_dret_i, csr_restore_dret_i };
  assign _0384_ = ~ { csr_save_cause_i, csr_save_cause_i };
  assign _0392_ = ~ { _3822_, _3822_, _3822_, _3822_ };
  assign _0394_ = ~ { _3822_, _3822_, _3822_, _3822_, _3822_, _3822_, _3822_, _3822_, _3822_, _3822_, _3822_, _3822_ };
  assign _0393_ = ~ { _3823_, _3823_ };
  assign _0395_ = ~ { _3822_, _3822_ };
  assign _0396_ = ~ { _3748_, _3748_ };
  assign _0397_ = ~ { _3746_, _3746_ };
  assign _0245_ = ~ _3823_;
  assign _0185_ = ~ _3832_;
  assign _0398_ = ~ { _3826_, _3826_, _3826_, _3826_, _3826_, _3826_, _3826_, _3826_, _3826_, _3826_, _3826_, _3826_, _3826_, _3826_, _3826_, _3826_, _3826_, _3826_, _3826_, _3826_, _3826_, _3826_, _3826_, _3826_, _3826_, _3826_, _3826_, _3826_, _3826_, _3826_, _3826_, _3826_ };
  assign _0399_ = ~ { _3830_, _3830_, _3830_, _3830_, _3830_, _3830_, _3830_, _3830_, _3830_, _3830_, _3830_, _3830_, _3830_, _3830_, _3830_, _3830_, _3830_, _3830_, _3830_, _3830_, _3830_, _3830_, _3830_, _3830_, _3830_, _3830_, _3830_, _3830_, _3830_, _3830_, _3830_, _3830_ };
  assign _0183_ = ~ _3833_;
  assign _0182_ = ~ _3834_;
  assign _0221_ = ~ _3835_;
  assign _0189_ = ~ _3836_;
  assign _0171_ = ~ _3822_;
  assign _0174_ = ~ _3837_;
  assign _0170_ = ~ _3839_;
  assign _0224_ = ~ _3840_;
  assign _0175_ = ~ _3841_;
  assign _0173_ = ~ _3842_;
  assign _0184_ = ~ _3843_;
  assign _0401_ = ~ { csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int };
  assign _0400_ = ~ csr_we_int;
  assign _0402_ = ~ { csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int };
  assign _0410_ = ~ { csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i };
  assign _0411_ = ~ { mstatus_q[1], mstatus_q[1] };
  assign _2069_ = { _3732_, _3732_, _3732_, _3732_, _3732_, _3732_, _3732_, _3732_, _3732_, _3732_, _3732_, _3732_, _3732_, _3732_, _3732_, _3732_, _3732_, _3732_, _3732_, _3732_, _3732_, _3732_, _3732_, _3732_, _3732_, _3732_, _3732_, _3732_, _3732_, _3732_, _3732_, _3732_ } | _0218_;
  assign _2072_ = { _0161_, _0161_, _0161_, _0161_, _0161_, _0161_, _0161_, _0161_, _0161_, _0161_, _0161_, _0161_, _0161_, _0161_, _0161_, _0161_, _0161_, _0161_, _0161_, _0161_, _0161_, _0161_, _0161_, _0161_, _0161_, _0161_, _0161_, _0161_, _0161_, _0161_, _0161_, _0161_ } | _0219_;
  assign _2101_ = _1998_ | _0225_;
  assign _2111_ = _0431_ | _0227_;
  assign _2138_ = { _0025_, _0025_, _0025_ } | _0236_;
  assign _2144_ = { _1998_, _1998_, _1998_ } | _0238_;
  assign _2153_ = { _2002_, _2002_, _2002_ } | _0241_;
  assign _2156_ = { _0435_, _0435_, _0435_ } | _0242_;
  assign _2159_ = { _0433_, _0433_, _0433_ } | _0243_;
  assign _2213_ = { _0441_, _0441_, _0441_ } | _0254_;
  assign _2228_ = { _2014_, _2014_, _2014_ } | _0258_;
  assign _2231_ = { _0443_, _0443_, _0443_ } | _0259_;
  assign _2234_ = { _0445_, _0445_, _0445_ } | _0260_;
  assign _2237_ = { _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_ } | _0261_;
  assign _2240_ = { _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_ } | _0262_;
  assign _2243_ = { _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_ } | _0263_;
  assign _2246_ = { _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_ } | _0264_;
  assign _2249_ = { _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_ } | _0265_;
  assign _2252_ = { _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_ } | _0266_;
  assign _2255_ = { _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_ } | _0267_;
  assign _2258_ = { _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_ } | _0268_;
  assign _2261_ = { _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_ } | _0269_;
  assign _2264_ = { _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_ } | _0270_;
  assign _2267_ = { _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_ } | _0271_;
  assign _2270_ = { _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_ } | _0272_;
  assign _2279_ = _3741_ | _0178_;
  assign _2280_ = _2008_ | _0273_;
  assign _2293_ = _0453_ | _0275_;
  assign _2307_ = _0455_ | _0277_;
  assign _2310_ = _0457_ | _0278_;
  assign _2313_ = _0459_ | _0279_;
  assign _2347_ = { _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_ } | _0280_;
  assign _2350_ = { _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_ } | _0281_;
  assign _2353_ = { _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_ } | _0282_;
  assign _2356_ = { _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_ } | _0283_;
  assign _2359_ = { _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_ } | _0284_;
  assign _2362_ = { _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_ } | _0285_;
  assign _2365_ = { _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_ } | _0286_;
  assign _2368_ = { _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_ } | _0287_;
  assign _2371_ = { _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_ } | _0288_;
  assign _2374_ = { _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_ } | _0289_;
  assign _2377_ = { _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_ } | _0290_;
  assign _2380_ = { _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_ } | _0291_;
  assign _2383_ = { _3743_, _3743_, _3743_, _3743_, _3743_, _3743_, _3743_, _3743_, _3743_ } | _0292_;
  assign _2386_ = { _3827_, _3827_, _3827_, _3827_, _3827_, _3827_, _3827_, _3827_, _3827_ } | _0293_;
  assign _2389_ = { _2022_, _2022_, _2022_, _2022_, _2022_, _2022_, _2022_, _2022_, _2022_ } | _0294_;
  assign _2392_ = { _3847_, _3847_, _3847_, _3847_, _3847_, _3847_, _3847_, _3847_, _3847_ } | _0295_;
  assign _2395_ = { _0031_, _0031_, _0031_, _0031_, _0031_, _0031_, _0031_, _0031_, _0031_ } | _0296_;
  assign _2398_ = { _0033_, _0033_, _0033_, _0033_, _0033_, _0033_, _0033_, _0033_, _0033_ } | _0297_;
  assign _2401_ = { _2018_, _2018_, _2018_, _2018_, _2018_, _2018_, _2018_, _2018_, _2018_ } | _0298_;
  assign _2404_ = { _0461_, _0461_, _0461_, _0461_, _0461_, _0461_, _0461_, _0461_, _0461_ } | _0299_;
  assign _2407_ = { _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_ } | _0300_;
  assign _2410_ = { _0045_, _0045_, _0045_, _0045_, _0045_, _0045_, _0045_, _0045_, _0045_ } | _0301_;
  assign _2413_ = { _0063_, _0063_, _0063_, _0063_, _0063_, _0063_, _0063_, _0063_, _0063_ } | _0302_;
  assign _2416_ = { _2020_, _2020_, _2020_, _2020_, _2020_, _2020_, _2020_, _2020_, _2020_ } | _0303_;
  assign _2419_ = { _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_ } | _0304_;
  assign _2422_ = { _3889_, _3889_, _3889_, _3889_, _3889_, _3889_, _3889_, _3889_, _3889_ } | _0305_;
  assign _2425_ = { _3891_, _3891_, _3891_, _3891_, _3891_, _3891_, _3891_, _3891_, _3891_ } | _0306_;
  assign _2428_ = { _2006_, _2006_, _2006_, _2006_, _2006_, _2006_, _2006_, _2006_, _2006_ } | _0307_;
  assign _2431_ = { _0463_, _0463_, _0463_, _0463_, _0463_, _0463_, _0463_, _0463_, _0463_ } | _0308_;
  assign _2434_ = { _0465_, _0465_, _0465_, _0465_, _0465_, _0465_, _0465_, _0465_, _0465_ } | _0309_;
  assign _2437_ = { _3827_, _3827_, _3827_ } | _0310_;
  assign _2441_ = { _3847_, _3847_, _3847_ } | _0311_;
  assign _2445_ = { _2018_, _2018_, _2018_ } | _0312_;
  assign _2448_ = { _0467_, _0467_, _0467_ } | _0313_;
  assign _2461_ = { _0469_, _0469_, _0469_ } | _0316_;
  assign _2464_ = { _0471_, _0471_, _0471_ } | _0317_;
  assign _2117_ = { _3743_, _3743_, _3743_ } | _0229_;
  assign _2123_ = { _1994_, _1994_, _1994_ } | _0231_;
  assign _2129_ = { _0031_, _0031_, _0031_ } | _0233_;
  assign _2132_ = { _1996_, _1996_, _1996_ } | _0234_;
  assign _2135_ = { _0429_, _0429_, _0429_ } | _0235_;
  assign _2475_ = { _3893_, _3893_, _3893_ } | _0318_;
  assign _2141_ = { _0045_, _0045_, _0045_ } | _0237_;
  assign _2479_ = { _2004_, _2004_, _2004_ } | _0319_;
  assign _2147_ = { _0053_, _0053_, _0053_ } | _0239_;
  assign _2487_ = { _2006_, _2006_, _2006_ } | _0321_;
  assign _2490_ = { _0437_, _0437_, _0437_ } | _0322_;
  assign _2493_ = { _0439_, _0439_, _0439_ } | _0323_;
  assign _2301_ = _2020_ | _0276_;
  assign _2510_ = _0473_ | _0324_;
  assign _2114_ = _0433_ | _0228_;
  assign _2078_ = _3831_ | _0187_;
  assign _2081_ = _1994_ | _0220_;
  assign _2089_ = _1996_ | _0222_;
  assign _2092_ = _0429_ | _0223_;
  assign _2172_ = _3893_ | _0180_;
  assign _2178_ = _2004_ | _0244_;
  assign _2187_ = _2006_ | _0246_;
  assign _2190_ = _0437_ | _0247_;
  assign _2193_ = _0439_ | _0248_;
  assign _2196_ = { _0021_, _0021_, _0021_ } | _0249_;
  assign _2530_ = { _3738_, _3738_, _3738_ } | _0325_;
  assign _2199_ = { _3741_, _3741_, _3741_ } | _0250_;
  assign _2202_ = { _2008_, _2008_, _2008_ } | _0251_;
  assign _2120_ = { _3831_, _3831_, _3831_ } | _0230_;
  assign _2206_ = { _0033_, _0033_, _0033_ } | _0252_;
  assign _2126_ = { _0041_, _0041_, _0041_ } | _0232_;
  assign _2210_ = { _2010_, _2010_, _2010_ } | _0253_;
  assign _2539_ = { _0475_, _0475_, _0475_ } | _0326_;
  assign _2216_ = { _0029_, _0029_, _0029_ } | _0255_;
  assign _2543_ = { _0039_, _0039_, _0039_ } | _0327_;
  assign _2219_ = { _0063_, _0063_, _0063_ } | _0256_;
  assign _2222_ = { _2012_, _2012_, _2012_ } | _0257_;
  assign _2454_ = { _3838_, _3838_, _3838_ } | _0314_;
  assign _2150_ = { _3889_, _3889_, _3889_ } | _0240_;
  assign _2484_ = { _3891_, _3891_, _3891_ } | _0320_;
  assign _2458_ = { _2000_, _2000_, _2000_ } | _0315_;
  assign _2552_ = { _0477_, _0477_, _0477_ } | _0328_;
  assign _2555_ = { _0479_, _0479_, _0479_ } | _0329_;
  assign _2075_ = _3743_ | _0179_;
  assign _2276_ = _3827_ | _0181_;
  assign _2559_ = _2024_ | _0330_;
  assign _2283_ = _3847_ | _0186_;
  assign _2290_ = _2018_ | _0274_;
  assign _2565_ = _0481_ | _0331_;
  assign _2570_ = _2012_ | _0332_;
  assign _2108_ = _2000_ | _0226_;
  assign _2576_ = _0469_ | _0333_;
  assign _2579_ = _0483_ | _0334_;
  assign _2583_ = _0157_ | _0335_;
  assign _2612_ = { nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0 } | _0364_;
  assign _2615_ = { nmi_mode_i_t0, nmi_mode_i_t0 } | _0365_;
  assign _2610_ = nmi_mode_i_t0 | _0363_;
  assign _2618_ = { csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0 } | _0366_;
  assign _2621_ = { csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0 } | _0367_;
  assign _2627_ = { nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0 } | _0369_;
  assign _2630_ = { debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0 } | _0370_;
  assign _2638_ = { debug_mode_i_t0, debug_mode_i_t0 } | _0373_;
  assign _2635_ = { debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0 } | _0372_;
  assign _2648_ = { debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0 } | _0376_;
  assign _2651_ = { debug_csr_save_i_t0, debug_csr_save_i_t0 } | _0377_;
  assign _2657_ = { debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0 } | _0378_;
  assign _2645_ = { debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0 } | _0375_;
  assign _2643_ = debug_csr_save_i_t0 | _0374_;
  assign _2663_ = { debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0 } | _0379_;
  assign _2666_ = { csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0 } | _0380_;
  assign _2669_ = { csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0 } | _0381_;
  assign _2672_ = { csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0 } | _0382_;
  assign _2624_ = { csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0 } | _0368_;
  assign _2689_ = { csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0 } | _0385_;
  assign _2692_ = { csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0 } | _0386_;
  assign _2695_ = { csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0 } | _0387_;
  assign _2701_ = { csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0 } | _0388_;
  assign _2704_ = { csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0 } | _0389_;
  assign _2676_ = { csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0 } | _0383_;
  assign _2601_ = csr_restore_mret_i_t0 | _0360_;
  assign _2604_ = csr_restore_dret_i_t0 | _0361_;
  assign _2607_ = csr_save_cause_i_t0 | _0362_;
  assign _2633_ = debug_mode_i_t0 | _0371_;
  assign _2710_ = { csr_restore_mret_i_t0, csr_restore_mret_i_t0 } | _0390_;
  assign _2713_ = { csr_restore_dret_i_t0, csr_restore_dret_i_t0 } | _0391_;
  assign _2681_ = { csr_save_cause_i_t0, csr_save_cause_i_t0 } | _0384_;
  assign _2717_ = { _0025_, _0025_, _0025_, _0025_ } | _0392_;
  assign _2725_ = { _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_ } | _0394_;
  assign _2720_ = { _0059_, _0059_ } | _0393_;
  assign _2729_ = { _0025_, _0025_ } | _0395_;
  assign _2734_ = { _3749_, _3749_ } | _0396_;
  assign _2737_ = { _3747_, _3747_ } | _0397_;
  assign _2184_ = _0059_ | _0245_;
  assign _2273_ = _0021_ | _0185_;
  assign _2740_ = { _3827_, _3827_, _3827_, _3827_, _3827_, _3827_, _3827_, _3827_, _3827_, _3827_, _3827_, _3827_, _3827_, _3827_, _3827_, _3827_, _3827_, _3827_, _3827_, _3827_, _3827_, _3827_, _3827_, _3827_, _3827_, _3827_, _3827_, _3827_, _3827_, _3827_, _3827_, _3827_ } | _0398_;
  assign _2743_ = { _3831_, _3831_, _3831_, _3831_, _3831_, _3831_, _3831_, _3831_, _3831_, _3831_, _3831_, _3831_, _3831_, _3831_, _3831_, _3831_, _3831_, _3831_, _3831_, _3831_, _3831_, _3831_, _3831_, _3831_, _3831_, _3831_, _3831_, _3831_, _3831_, _3831_, _3831_, _3831_ } | _0399_;
  assign _2084_ = _0041_ | _0183_;
  assign _2287_ = _0033_ | _0182_;
  assign _2086_ = _0031_ | _0221_;
  assign _2166_ = _0029_ | _0189_;
  assign _2095_ = _0025_ | _0171_;
  assign _2104_ = _3838_ | _0174_;
  assign _2298_ = _0063_ | _0170_;
  assign _2098_ = _0039_ | _0224_;
  assign _2175_ = _0045_ | _0175_;
  assign _2181_ = _0053_ | _0173_;
  assign _2506_ = _0051_ | _0184_;
  assign _2748_ = { csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0 } | _0401_;
  assign _2746_ = csr_we_int_t0 | _0400_;
  assign _2754_ = { csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0 } | _0402_;
  assign _2757_ = { csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0 } | _0410_;
  assign _2760_ = { mstatus_q_t0[1], mstatus_q_t0[1] } | _0411_;
  assign _2070_ = { _3732_, _3732_, _3732_, _3732_, _3732_, _3732_, _3732_, _3732_, _3732_, _3732_, _3732_, _3732_, _3732_, _3732_, _3732_, _3732_, _3732_, _3732_, _3732_, _3732_, _3732_, _3732_, _3732_, _3732_, _3732_, _3732_, _3732_, _3732_, _3732_, _3732_, _3732_, _3732_ } | { _3731_, _3731_, _3731_, _3731_, _3731_, _3731_, _3731_, _3731_, _3731_, _3731_, _3731_, _3731_, _3731_, _3731_, _3731_, _3731_, _3731_, _3731_, _3731_, _3731_, _3731_, _3731_, _3731_, _3731_, _3731_, _3731_, _3731_, _3731_, _3731_, _3731_, _3731_, _3731_ };
  assign _2073_ = { _0161_, _0161_, _0161_, _0161_, _0161_, _0161_, _0161_, _0161_, _0161_, _0161_, _0161_, _0161_, _0161_, _0161_, _0161_, _0161_, _0161_, _0161_, _0161_, _0161_, _0161_, _0161_, _0161_, _0161_, _0161_, _0161_, _0161_, _0161_, _0161_, _0161_, _0161_, _0161_ } | { _0160_, _0160_, _0160_, _0160_, _0160_, _0160_, _0160_, _0160_, _0160_, _0160_, _0160_, _0160_, _0160_, _0160_, _0160_, _0160_, _0160_, _0160_, _0160_, _0160_, _0160_, _0160_, _0160_, _0160_, _0160_, _0160_, _0160_, _0160_, _0160_, _0160_, _0160_, _0160_ };
  assign _2102_ = _1998_ | _1997_;
  assign _2112_ = _0431_ | _0430_;
  assign _2139_ = { _0025_, _0025_, _0025_ } | { _3822_, _3822_, _3822_ };
  assign _2145_ = { _1998_, _1998_, _1998_ } | { _1997_, _1997_, _1997_ };
  assign _2154_ = { _2002_, _2002_, _2002_ } | { _2001_, _2001_, _2001_ };
  assign _2157_ = { _0435_, _0435_, _0435_ } | { _0434_, _0434_, _0434_ };
  assign _2160_ = { _0433_, _0433_, _0433_ } | { _0432_, _0432_, _0432_ };
  assign _2214_ = { _0441_, _0441_, _0441_ } | { _0440_, _0440_, _0440_ };
  assign _2229_ = { _2014_, _2014_, _2014_ } | { _2013_, _2013_, _2013_ };
  assign _2232_ = { _0443_, _0443_, _0443_ } | { _0442_, _0442_, _0442_ };
  assign _2235_ = { _0445_, _0445_, _0445_ } | { _0444_, _0444_, _0444_ };
  assign _2238_ = { _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_ } | { _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_ };
  assign _2241_ = { _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_ } | { _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_ };
  assign _2244_ = { _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_ } | { _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_ };
  assign _2247_ = { _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_ } | { _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_ };
  assign _2250_ = { _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_ } | { _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_ };
  assign _2253_ = { _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_ } | { _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_ };
  assign _2256_ = { _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_ } | { _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_ };
  assign _2259_ = { _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_ } | { _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_ };
  assign _2262_ = { _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_ } | { _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_ };
  assign _2265_ = { _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_ } | { _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_ };
  assign _2268_ = { _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_ } | { _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_ };
  assign _2271_ = { _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_ } | { _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_ };
  assign _2281_ = _2008_ | _2007_;
  assign _2294_ = _0453_ | _0452_;
  assign _2308_ = _0455_ | _0454_;
  assign _2311_ = _0457_ | _0456_;
  assign _2314_ = _0459_ | _0458_;
  assign _2348_ = { _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_ } | { _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_, _3932_ };
  assign _2351_ = { _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_ } | { _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_ };
  assign _2354_ = { _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_ } | { _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_, _3938_ };
  assign _2357_ = { _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_ } | { _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_, _3936_ };
  assign _2360_ = { _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_ } | { _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_ };
  assign _2363_ = { _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_ } | { _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_, _3944_ };
  assign _2366_ = { _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_ } | { _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_, _3942_ };
  assign _2369_ = { _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_ } | { _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_, _3948_ };
  assign _2372_ = { _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_ } | { _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_, _3952_ };
  assign _2375_ = { _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_ } | { _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_, _2015_ };
  assign _2378_ = { _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_ } | { _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_, _0448_ };
  assign _2381_ = { _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_ } | { _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_, _0450_ };
  assign _2384_ = { _3743_, _3743_, _3743_, _3743_, _3743_, _3743_, _3743_, _3743_, _3743_ } | { _3742_, _3742_, _3742_, _3742_, _3742_, _3742_, _3742_, _3742_, _3742_ };
  assign _2387_ = { _3827_, _3827_, _3827_, _3827_, _3827_, _3827_, _3827_, _3827_, _3827_ } | { _3826_, _3826_, _3826_, _3826_, _3826_, _3826_, _3826_, _3826_, _3826_ };
  assign _2390_ = { _2022_, _2022_, _2022_, _2022_, _2022_, _2022_, _2022_, _2022_, _2022_ } | { _2021_, _2021_, _2021_, _2021_, _2021_, _2021_, _2021_, _2021_, _2021_ };
  assign _2393_ = { _3847_, _3847_, _3847_, _3847_, _3847_, _3847_, _3847_, _3847_, _3847_ } | { _3846_, _3846_, _3846_, _3846_, _3846_, _3846_, _3846_, _3846_, _3846_ };
  assign _2396_ = { _0031_, _0031_, _0031_, _0031_, _0031_, _0031_, _0031_, _0031_, _0031_ } | { _3835_, _3835_, _3835_, _3835_, _3835_, _3835_, _3835_, _3835_, _3835_ };
  assign _2399_ = { _0033_, _0033_, _0033_, _0033_, _0033_, _0033_, _0033_, _0033_, _0033_ } | { _3834_, _3834_, _3834_, _3834_, _3834_, _3834_, _3834_, _3834_, _3834_ };
  assign _2402_ = { _2018_, _2018_, _2018_, _2018_, _2018_, _2018_, _2018_, _2018_, _2018_ } | { _2017_, _2017_, _2017_, _2017_, _2017_, _2017_, _2017_, _2017_, _2017_ };
  assign _2405_ = { _0461_, _0461_, _0461_, _0461_, _0461_, _0461_, _0461_, _0461_, _0461_ } | { _0460_, _0460_, _0460_, _0460_, _0460_, _0460_, _0460_, _0460_, _0460_ };
  assign _2408_ = { _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_ } | { _3822_, _3822_, _3822_, _3822_, _3822_, _3822_, _3822_, _3822_, _3822_ };
  assign _2411_ = { _0045_, _0045_, _0045_, _0045_, _0045_, _0045_, _0045_, _0045_, _0045_ } | { _3841_, _3841_, _3841_, _3841_, _3841_, _3841_, _3841_, _3841_, _3841_ };
  assign _2414_ = { _0063_, _0063_, _0063_, _0063_, _0063_, _0063_, _0063_, _0063_, _0063_ } | { _3839_, _3839_, _3839_, _3839_, _3839_, _3839_, _3839_, _3839_, _3839_ };
  assign _2417_ = { _2020_, _2020_, _2020_, _2020_, _2020_, _2020_, _2020_, _2020_, _2020_ } | { _2019_, _2019_, _2019_, _2019_, _2019_, _2019_, _2019_, _2019_, _2019_ };
  assign _2420_ = { _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_ } | { _3842_, _3842_, _3842_, _3842_, _3842_, _3842_, _3842_, _3842_, _3842_ };
  assign _2423_ = { _3889_, _3889_, _3889_, _3889_, _3889_, _3889_, _3889_, _3889_, _3889_ } | { _3888_, _3888_, _3888_, _3888_, _3888_, _3888_, _3888_, _3888_, _3888_ };
  assign _2426_ = { _3891_, _3891_, _3891_, _3891_, _3891_, _3891_, _3891_, _3891_, _3891_ } | { _3890_, _3890_, _3890_, _3890_, _3890_, _3890_, _3890_, _3890_, _3890_ };
  assign _2429_ = { _2006_, _2006_, _2006_, _2006_, _2006_, _2006_, _2006_, _2006_, _2006_ } | { _2005_, _2005_, _2005_, _2005_, _2005_, _2005_, _2005_, _2005_, _2005_ };
  assign _2432_ = { _0463_, _0463_, _0463_, _0463_, _0463_, _0463_, _0463_, _0463_, _0463_ } | { _0462_, _0462_, _0462_, _0462_, _0462_, _0462_, _0462_, _0462_, _0462_ };
  assign _2435_ = { _0465_, _0465_, _0465_, _0465_, _0465_, _0465_, _0465_, _0465_, _0465_ } | { _0464_, _0464_, _0464_, _0464_, _0464_, _0464_, _0464_, _0464_, _0464_ };
  assign _2438_ = { _3827_, _3827_, _3827_ } | { _3826_, _3826_, _3826_ };
  assign _2442_ = { _3847_, _3847_, _3847_ } | { _3846_, _3846_, _3846_ };
  assign _2446_ = { _2018_, _2018_, _2018_ } | { _2017_, _2017_, _2017_ };
  assign _2449_ = { _0467_, _0467_, _0467_ } | { _0466_, _0466_, _0466_ };
  assign _2462_ = { _0469_, _0469_, _0469_ } | { _0468_, _0468_, _0468_ };
  assign _2465_ = { _0471_, _0471_, _0471_ } | { _0470_, _0470_, _0470_ };
  assign _2118_ = { _3743_, _3743_, _3743_ } | { _3742_, _3742_, _3742_ };
  assign _2124_ = { _1994_, _1994_, _1994_ } | { _1993_, _1993_, _1993_ };
  assign _2130_ = { _0031_, _0031_, _0031_ } | { _3835_, _3835_, _3835_ };
  assign _2133_ = { _1996_, _1996_, _1996_ } | { _1995_, _1995_, _1995_ };
  assign _2136_ = { _0429_, _0429_, _0429_ } | { _0428_, _0428_, _0428_ };
  assign _2476_ = { _3893_, _3893_, _3893_ } | { _3892_, _3892_, _3892_ };
  assign _2142_ = { _0045_, _0045_, _0045_ } | { _3841_, _3841_, _3841_ };
  assign _2480_ = { _2004_, _2004_, _2004_ } | { _2003_, _2003_, _2003_ };
  assign _2148_ = { _0053_, _0053_, _0053_ } | { _3842_, _3842_, _3842_ };
  assign _2488_ = { _2006_, _2006_, _2006_ } | { _2005_, _2005_, _2005_ };
  assign _2491_ = { _0437_, _0437_, _0437_ } | { _0436_, _0436_, _0436_ };
  assign _2494_ = { _0439_, _0439_, _0439_ } | { _0438_, _0438_, _0438_ };
  assign _2302_ = _2020_ | _2019_;
  assign _2511_ = _0473_ | _0472_;
  assign _2115_ = _0433_ | _0432_;
  assign _2079_ = _3831_ | _3830_;
  assign _2082_ = _1994_ | _1993_;
  assign _2090_ = _1996_ | _1995_;
  assign _2093_ = _0429_ | _0428_;
  assign _2173_ = _3893_ | _3892_;
  assign _2179_ = _2004_ | _2003_;
  assign _2188_ = _2006_ | _2005_;
  assign _2191_ = _0437_ | _0436_;
  assign _2194_ = _0439_ | _0438_;
  assign _2197_ = { _0021_, _0021_, _0021_ } | { _3832_, _3832_, _3832_ };
  assign _2531_ = { _3738_, _3738_, _3738_ } | { _3737_, _3737_, _3737_ };
  assign _2200_ = { _3741_, _3741_, _3741_ } | { _3740_, _3740_, _3740_ };
  assign _2203_ = { _2008_, _2008_, _2008_ } | { _2007_, _2007_, _2007_ };
  assign _2121_ = { _3831_, _3831_, _3831_ } | { _3830_, _3830_, _3830_ };
  assign _2207_ = { _0033_, _0033_, _0033_ } | { _3834_, _3834_, _3834_ };
  assign _2127_ = { _0041_, _0041_, _0041_ } | { _3833_, _3833_, _3833_ };
  assign _2211_ = { _2010_, _2010_, _2010_ } | { _2009_, _2009_, _2009_ };
  assign _2540_ = { _0475_, _0475_, _0475_ } | { _0474_, _0474_, _0474_ };
  assign _2217_ = { _0029_, _0029_, _0029_ } | { _3836_, _3836_, _3836_ };
  assign _2544_ = { _0039_, _0039_, _0039_ } | { _3840_, _3840_, _3840_ };
  assign _2220_ = { _0063_, _0063_, _0063_ } | { _3839_, _3839_, _3839_ };
  assign _2223_ = { _2012_, _2012_, _2012_ } | { _2011_, _2011_, _2011_ };
  assign _2455_ = { _3838_, _3838_, _3838_ } | { _3837_, _3837_, _3837_ };
  assign _2151_ = { _3889_, _3889_, _3889_ } | { _3888_, _3888_, _3888_ };
  assign _2485_ = { _3891_, _3891_, _3891_ } | { _3890_, _3890_, _3890_ };
  assign _2459_ = { _2000_, _2000_, _2000_ } | { _1999_, _1999_, _1999_ };
  assign _2553_ = { _0477_, _0477_, _0477_ } | { _0476_, _0476_, _0476_ };
  assign _2556_ = { _0479_, _0479_, _0479_ } | { _0478_, _0478_, _0478_ };
  assign _2076_ = _3743_ | _3742_;
  assign _2277_ = _3827_ | _3826_;
  assign _2560_ = _2024_ | _2023_;
  assign _2284_ = _3847_ | _3846_;
  assign _2291_ = _2018_ | _2017_;
  assign _2566_ = _0481_ | _0480_;
  assign _2571_ = _2012_ | _2011_;
  assign _2107_ = _3889_ | _3888_;
  assign _2109_ = _2000_ | _1999_;
  assign _2577_ = _0469_ | _0468_;
  assign _2580_ = _0483_ | _0482_;
  assign _2582_ = _0159_ | _0158_;
  assign _2613_ = { nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0 } | { nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i };
  assign _2616_ = { nmi_mode_i_t0, nmi_mode_i_t0 } | { nmi_mode_i, nmi_mode_i };
  assign _2611_ = nmi_mode_i_t0 | nmi_mode_i;
  assign _2619_ = { csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0 } | { csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i };
  assign _2622_ = { csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0 } | { csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i };
  assign _2628_ = { nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0 } | { nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i };
  assign _2631_ = { debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0 } | { debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i };
  assign _2639_ = { debug_mode_i_t0, debug_mode_i_t0 } | { debug_mode_i, debug_mode_i };
  assign _2636_ = { debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0 } | { debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i };
  assign _2649_ = { debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0 } | { debug_csr_save_i, debug_csr_save_i, debug_csr_save_i };
  assign _2652_ = { debug_csr_save_i_t0, debug_csr_save_i_t0 } | { debug_csr_save_i, debug_csr_save_i };
  assign _2658_ = { debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0 } | { debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i };
  assign _2646_ = { debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0 } | { debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i };
  assign _2644_ = debug_csr_save_i_t0 | debug_csr_save_i;
  assign _2664_ = { debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0 } | { debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i };
  assign _2667_ = { csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0 } | { csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i };
  assign _2670_ = { csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0 } | { csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i };
  assign _2673_ = { csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0 } | { csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i };
  assign _2625_ = { csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0 } | { csr_save_cause_i, csr_save_cause_i, csr_save_cause_i };
  assign _2690_ = { csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0 } | { csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i };
  assign _2693_ = { csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0 } | { csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i };
  assign _2696_ = { csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0 } | { csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i };
  assign _2702_ = { csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0 } | { csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i };
  assign _2705_ = { csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0 } | { csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i };
  assign _2677_ = { csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0 } | { csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i };
  assign _2602_ = csr_restore_mret_i_t0 | csr_restore_mret_i;
  assign _2605_ = csr_restore_dret_i_t0 | csr_restore_dret_i;
  assign _2608_ = csr_save_cause_i_t0 | csr_save_cause_i;
  assign _2634_ = debug_mode_i_t0 | debug_mode_i;
  assign _2711_ = { csr_restore_mret_i_t0, csr_restore_mret_i_t0 } | { csr_restore_mret_i, csr_restore_mret_i };
  assign _2714_ = { csr_restore_dret_i_t0, csr_restore_dret_i_t0 } | { csr_restore_dret_i, csr_restore_dret_i };
  assign _2682_ = { csr_save_cause_i_t0, csr_save_cause_i_t0 } | { csr_save_cause_i, csr_save_cause_i };
  assign _2718_ = { _0025_, _0025_, _0025_, _0025_ } | { _3822_, _3822_, _3822_, _3822_ };
  assign _2726_ = { _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_ } | { _3822_, _3822_, _3822_, _3822_, _3822_, _3822_, _3822_, _3822_, _3822_, _3822_, _3822_, _3822_ };
  assign _2721_ = { _0059_, _0059_ } | { _3823_, _3823_ };
  assign _2730_ = { _0025_, _0025_ } | { _3822_, _3822_ };
  assign _2735_ = { _3749_, _3749_ } | { _3748_, _3748_ };
  assign _2738_ = { _3747_, _3747_ } | { _3746_, _3746_ };
  assign _2185_ = _0059_ | _3823_;
  assign _2274_ = _0021_ | _3832_;
  assign _2741_ = { _3827_, _3827_, _3827_, _3827_, _3827_, _3827_, _3827_, _3827_, _3827_, _3827_, _3827_, _3827_, _3827_, _3827_, _3827_, _3827_, _3827_, _3827_, _3827_, _3827_, _3827_, _3827_, _3827_, _3827_, _3827_, _3827_, _3827_, _3827_, _3827_, _3827_, _3827_, _3827_ } | { _3826_, _3826_, _3826_, _3826_, _3826_, _3826_, _3826_, _3826_, _3826_, _3826_, _3826_, _3826_, _3826_, _3826_, _3826_, _3826_, _3826_, _3826_, _3826_, _3826_, _3826_, _3826_, _3826_, _3826_, _3826_, _3826_, _3826_, _3826_, _3826_, _3826_, _3826_, _3826_ };
  assign _2744_ = { _3831_, _3831_, _3831_, _3831_, _3831_, _3831_, _3831_, _3831_, _3831_, _3831_, _3831_, _3831_, _3831_, _3831_, _3831_, _3831_, _3831_, _3831_, _3831_, _3831_, _3831_, _3831_, _3831_, _3831_, _3831_, _3831_, _3831_, _3831_, _3831_, _3831_, _3831_, _3831_ } | { _3830_, _3830_, _3830_, _3830_, _3830_, _3830_, _3830_, _3830_, _3830_, _3830_, _3830_, _3830_, _3830_, _3830_, _3830_, _3830_, _3830_, _3830_, _3830_, _3830_, _3830_, _3830_, _3830_, _3830_, _3830_, _3830_, _3830_, _3830_, _3830_, _3830_, _3830_, _3830_ };
  assign _2085_ = _0041_ | _3833_;
  assign _2288_ = _0033_ | _3834_;
  assign _2087_ = _0031_ | _3835_;
  assign _2167_ = _0029_ | _3836_;
  assign _2096_ = _0025_ | _3822_;
  assign _2105_ = _3838_ | _3837_;
  assign _2299_ = _0063_ | _3839_;
  assign _2099_ = _0039_ | _3840_;
  assign _2176_ = _0045_ | _3841_;
  assign _2182_ = _0053_ | _3842_;
  assign _2507_ = _0051_ | _3843_;
  assign _2749_ = { csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0 } | { csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int };
  assign _2747_ = csr_we_int_t0 | csr_we_int;
  assign _2755_ = { csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0 } | { csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int };
  assign _2758_ = { csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0 } | { csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i };
  assign _2761_ = { mstatus_q_t0[1], mstatus_q_t0[1] } | { mstatus_q[1], mstatus_q[1] };
  assign _2763_ = _3751_ | _3750_;
  assign _0725_ = _3781_ & _2069_;
  assign _0728_ = _3242_ & _2072_;
  assign _0731_ = _0017_[63] & _2075_;
  assign _0734_ = _0019_[31] & _2078_;
  assign _0737_ = _3246_ & _2081_;
  assign _0740_ = dscratch1_q_t0[31] & _2084_;
  assign _0742_ = csr_depc_o_t0[31] & _2086_;
  assign _0745_ = _3252_ & _2089_;
  assign _0748_ = _3254_ & _2092_;
  assign _0751_ = mtval_q_t0[31] & _2095_;
  assign _0754_ = csr_mepc_o_t0[31] & _2098_;
  assign _0757_ = _3260_ & _2101_;
  assign _0760_ = mscratch_q_t0[31] & _2104_;
  assign _0765_ = _3266_ & _2108_;
  assign _0768_ = _3268_ & _2111_;
  assign _0771_ = _3270_ & _2114_;
  assign _0774_ = _0017_[42:40] & _2117_;
  assign _0777_ = _0019_[10:8] & _2120_;
  assign _0780_ = _3274_ & _2123_;
  assign _0783_ = dscratch1_q_t0[10:8] & _2126_;
  assign _0786_ = csr_depc_o_t0[10:8] & _2129_;
  assign _0789_ = _3280_ & _2132_;
  assign _0792_ = _3282_ & _2135_;
  assign _0795_ = mtval_q_t0[10:8] & _2138_;
  assign _0798_ = csr_mtvec_o_t0[10:8] & _2141_;
  assign _0801_ = _3288_ & _2144_;
  assign _0804_ = 3'h0 & _2147_;
  assign _0810_ = _3294_ & _2153_;
  assign _0813_ = _3296_ & _2156_;
  assign _0816_ = _3298_ & _2159_;
  assign _0819_ = _0017_[39] & _2075_;
  assign _0822_ = _0019_[7] & _2078_;
  assign _0825_ = _3302_ & _2081_;
  assign _0828_ = dscratch1_q_t0[7] & _2084_;
  assign _0831_ = dcsr_q_t0[7] & _2166_;
  assign _0834_ = _3308_ & _2086_;
  assign _0837_ = _3310_ & _2089_;
  assign _0840_ = _3312_ & _2092_;
  assign _0843_ = mtval_q_t0[7] & _2172_;
  assign _0846_ = csr_mtvec_o_t0[7] & _2175_;
  assign _0849_ = _3318_ & _2178_;
  assign _0852_ = mie_q_t0[16] & _2181_;
  assign _0857_ = _3324_ & _2184_;
  assign _0860_ = _3326_ & _2187_;
  assign _0863_ = _3328_ & _2190_;
  assign _0866_ = _3330_ & _2193_;
  assign _0869_ = \gen_trigger_regs.selected_tmatch_value_t0 [6:4] & _2196_;
  assign _0872_ = _0017_[38:36] & _2199_;
  assign _0875_ = _3334_ & _2202_;
  assign _0878_ = _0019_[6:4] & _2120_;
  assign _0881_ = dscratch0_q_t0[6:4] & _2206_;
  assign _0884_ = _3340_ & _2126_;
  assign _0887_ = _3342_ & _2210_;
  assign _0890_ = _3344_ & _2213_;
  assign _0893_ = dcsr_q_t0[6:4] & _2216_;
  assign _0896_ = { 2'h0, mcause_q_t0[4] } & _2219_;
  assign _0899_ = _3350_ & _2222_;
  assign _0902_ = csr_mtvec_o_t0[6:4] & _2141_;
  assign _0907_ = _3356_ & _2147_;
  assign _0910_ = _3358_ & _2228_;
  assign _0913_ = _3360_ & _2231_;
  assign _0916_ = _3362_ & _2234_;
  assign _0919_ = 32'd0 & _2237_;
  assign _0922_ = _3363_ & _2240_;
  assign _0925_ = 32'd0 & _2243_;
  assign _0928_ = _3367_ & _2246_;
  assign _0931_ = _3369_ & _2249_;
  assign _0934_ = 32'd0 & _2252_;
  assign _0937_ = _3373_ & _2255_;
  assign _0940_ = 32'd0 & _2258_;
  assign _0943_ = 32'd0 & _2261_;
  assign _0946_ = _3379_ & _2264_;
  assign _0949_ = _3381_ & _2267_;
  assign _0952_ = _3383_ & _2270_;
  assign _0955_ = \gen_trigger_regs.selected_tmatch_value_t0 [3] & _2273_;
  assign _0958_ = _0017_[3] & _2276_;
  assign _0961_ = _3387_ & _2279_;
  assign _0963_ = _3389_ & _2280_;
  assign _0966_ = mcountinhibit_t0[3] & _2283_;
  assign _0969_ = csr_depc_o_t0[3] & _2086_;
  assign _0972_ = _3395_ & _2287_;
  assign _0975_ = _3397_ & _2290_;
  assign _0978_ = _3399_ & _2293_;
  assign _0981_ = irq_software_i_t0 & _2095_;
  assign _0984_ = csr_mepc_o_t0[3] & _2098_;
  assign _0987_ = _3405_ & _2298_;
  assign _0990_ = _3407_ & _2301_;
  assign _0993_ = mie_q_t0[17] & _2181_;
  assign _0996_ = _3411_ & _2104_;
  assign _1001_ = _3415_ & _2184_;
  assign _1004_ = _3417_ & _2307_;
  assign _1007_ = _3419_ & _2310_;
  assign _1010_ = _3421_ & _2313_;
  assign _1013_ = _0017_[43] & _2075_;
  assign _1016_ = _0019_[11] & _2078_;
  assign _1019_ = _3425_ & _2081_;
  assign _1022_ = dscratch1_q_t0[11] & _2084_;
  assign _1025_ = dcsr_q_t0[11] & _2166_;
  assign _1028_ = _3431_ & _2086_;
  assign _1031_ = _3433_ & _2089_;
  assign _1034_ = _3435_ & _2092_;
  assign _1037_ = mtval_q_t0[11] & _2172_;
  assign _1040_ = csr_mtvec_o_t0[11] & _2175_;
  assign _1043_ = _3441_ & _2178_;
  assign _1046_ = mie_q_t0[15] & _2181_;
  assign _1051_ = _3447_ & _2184_;
  assign _1054_ = _3449_ & _2187_;
  assign _1057_ = _3451_ & _2190_;
  assign _1060_ = _3453_ & _2193_;
  assign _1063_ = _0017_[53] & _2075_;
  assign _1066_ = _0019_[21] & _2078_;
  assign _1069_ = _3457_ & _2081_;
  assign _1072_ = dscratch1_q_t0[21] & _2084_;
  assign _1074_ = dcsr_q_t0[21] & _2166_;
  assign _1077_ = _3463_ & _2086_;
  assign _1080_ = _3465_ & _2089_;
  assign _1083_ = _3467_ & _2092_;
  assign _1086_ = mtval_q_t0[21] & _2172_;
  assign _1089_ = csr_mtvec_o_t0[21] & _2175_;
  assign _1092_ = _3473_ & _2178_;
  assign _1095_ = mie_q_t0[5] & _2181_;
  assign _1100_ = _3479_ & _2184_;
  assign _1103_ = _3481_ & _2187_;
  assign _1106_ = _3483_ & _2190_;
  assign _1109_ = _3485_ & _2193_;
  assign _1112_ = \mhpmcounter[11]_t0  & _2347_;
  assign _1115_ = _3486_ & _2350_;
  assign _1118_ = \mhpmcounter[8]_t0  & _2353_;
  assign _1121_ = _3490_ & _2356_;
  assign _1124_ = _3492_ & _2359_;
  assign _1127_ = \mhpmcounter[5]_t0  & _2362_;
  assign _1130_ = _3496_ & _2365_;
  assign _1133_ = \mhpmcounter[3]_t0  & _2368_;
  assign _1136_ = \mhpmcounter[0]_t0  & _2371_;
  assign _1139_ = _3502_ & _2374_;
  assign _1142_ = _3504_ & _2377_;
  assign _1145_ = _3506_ & _2380_;
  assign _1148_ = 9'h000 & _2383_;
  assign _1151_ = _0017_[30:22] & _2386_;
  assign _1154_ = _3510_ & _2389_;
  assign _1157_ = 9'h000 & _2392_;
  assign _1160_ = csr_depc_o_t0[30:22] & _2395_;
  assign _1163_ = _3516_ & _2398_;
  assign _1166_ = _3518_ & _2401_;
  assign _1169_ = _3520_ & _2404_;
  assign _1172_ = irq_fast_i_t0[14:6] & _2407_;
  assign _1175_ = csr_mtvec_o_t0[30:22] & _2410_;
  assign _1178_ = _3526_ & _2413_;
  assign _1181_ = _3528_ & _2416_;
  assign _1184_ = mie_q_t0[14:6] & _2419_;
  assign _1187_ = 9'h000 & _2422_;
  assign _1190_ = _3534_ & _2425_;
  assign _1193_ = _3536_ & _2428_;
  assign _1196_ = _3538_ & _2431_;
  assign _1199_ = _3540_ & _2434_;
  assign _1202_ = _0017_[15:13] & _2437_;
  assign _1205_ = _3542_ & _2117_;
  assign _1208_ = 3'h0 & _2441_;
  assign _1211_ = dscratch0_q_t0[15:13] & _2206_;
  assign _1214_ = _3548_ & _2445_;
  assign _1217_ = _3550_ & _2448_;
  assign _1220_ = dcsr_q_t0[15:13] & _2216_;
  assign _1223_ = csr_mepc_o_t0[15:13] & _2219_;
  assign _1226_ = _3556_ & _2222_;
  assign _1229_ = mscratch_q_t0[15:13] & _2454_;
  assign _1234_ = _3562_ & _2458_;
  assign _1237_ = _3564_ & _2461_;
  assign _1240_ = _3566_ & _2464_;
  assign _1243_ = _0017_[52:50] & _2117_;
  assign _1246_ = _0019_[20:18] & _2120_;
  assign _1249_ = _3570_ & _2123_;
  assign _1252_ = dscratch1_q_t0[20:18] & _2126_;
  assign _1255_ = dcsr_q_t0[20:18] & _2216_;
  assign _1258_ = _3576_ & _2129_;
  assign _1261_ = _3578_ & _2132_;
  assign _1264_ = _3580_ & _2135_;
  assign _1267_ = mtval_q_t0[20:18] & _2475_;
  assign _1270_ = csr_mtvec_o_t0[20:18] & _2141_;
  assign _1273_ = _3586_ & _2479_;
  assign _1276_ = mie_q_t0[4:2] & _2147_;
  assign _1281_ = _3592_ & _2484_;
  assign _1284_ = _3594_ & _2487_;
  assign _1287_ = _3596_ & _2490_;
  assign _1290_ = _3598_ & _2493_;
  assign _1293_ = _0017_[48] & _2075_;
  assign _1296_ = _0019_[16] & _2078_;
  assign _1299_ = _3602_ & _2081_;
  assign _1302_ = dscratch1_q_t0[16] & _2084_;
  assign _1304_ = csr_depc_o_t0[16] & _2086_;
  assign _1307_ = _3608_ & _2089_;
  assign _1310_ = _3610_ & _2092_;
  assign _1313_ = irq_fast_i_t0[0] & _2095_;
  assign _1316_ = csr_mepc_o_t0[16] & _2298_;
  assign _1319_ = _3616_ & _2301_;
  assign _1322_ = mscratch_q_t0[16] & _2104_;
  assign _1327_ = _3622_ & _2506_;
  assign _1330_ = _3624_ & _2108_;
  assign _1333_ = _3626_ & _2510_;
  assign _1336_ = _3628_ & _2114_;
  assign _1339_ = _0017_[49] & _2075_;
  assign _1342_ = _0019_[17] & _2078_;
  assign _1345_ = _3632_ & _2081_;
  assign _1348_ = dscratch1_q_t0[17] & _2084_;
  assign _1350_ = dcsr_q_t0[17] & _2166_;
  assign _1353_ = _3638_ & _2086_;
  assign _1356_ = _3640_ & _2089_;
  assign _1359_ = _3642_ & _2092_;
  assign _1362_ = mtval_q_t0[17] & _2172_;
  assign _1365_ = csr_mtvec_o_t0[17] & _2175_;
  assign _1368_ = _3648_ & _2178_;
  assign _1371_ = mie_q_t0[1] & _2181_;
  assign _1376_ = _3654_ & _2184_;
  assign _1379_ = _3656_ & _2187_;
  assign _1382_ = _3658_ & _2190_;
  assign _1385_ = _3660_ & _2193_;
  assign _1388_ = \gen_trigger_regs.selected_tmatch_value_t0 [2:0] & _2196_;
  assign _1391_ = _0017_[34:32] & _2530_;
  assign _1394_ = _3664_ & _2199_;
  assign _1397_ = _3666_ & _2202_;
  assign _1400_ = _0019_[2:0] & _2120_;
  assign _1403_ = dscratch0_q_t0[2:0] & _2206_;
  assign _1406_ = _3672_ & _2126_;
  assign _1409_ = _3674_ & _2210_;
  assign _1412_ = _3676_ & _2539_;
  assign _1415_ = dcsr_q_t0[2:0] & _2216_;
  assign _1418_ = csr_mepc_o_t0[2:0] & _2543_;
  assign _1421_ = _3682_ & _2219_;
  assign _1424_ = _3684_ & _2222_;
  assign _1427_ = mscratch_q_t0[2:0] & _2454_;
  assign _0807_ = 3'h0 & _2150_;
  assign _1432_ = _3690_ & _2484_;
  assign _1434_ = _3692_ & _2458_;
  assign _1437_ = _3694_ & _2552_;
  assign _1440_ = _3696_ & _2555_;
  assign _1445_ = _0017_[12] & _2276_;
  assign _1448_ = _3700_ & _2559_;
  assign _1451_ = mcountinhibit_t0[12] & _2283_;
  assign _1454_ = dscratch0_q_t0[12] & _2287_;
  assign _1457_ = _3706_ & _2290_;
  assign _1460_ = _3708_ & _2565_;
  assign _1463_ = dcsr_q_t0[12] & _2166_;
  assign _1466_ = csr_mepc_o_t0[12] & _2298_;
  assign _1469_ = _3714_ & _2570_;
  assign _1472_ = mscratch_q_t0[12] & _2104_;
  assign _1477_ = _3720_ & _2184_;
  assign _1480_ = _3722_ & _2108_;
  assign _1483_ = _3724_ & _2576_;
  assign _1486_ = _3726_ & _2579_;
  assign _1491_ = _3727_ & _2583_;
  assign _1537_ = _0011_[5] & _2601_;
  assign _1540_ = _3787_ & _2604_;
  assign _1543_ = _3789_ & _2607_;
  assign _1546_ = _0007_ & _2610_;
  assign _1548_ = { csr_wdata_int_t0[31:1], 1'h0 } & _2612_;
  assign _1551_ = _0009_ & _2610_;
  assign _1553_ = 2'h0 & _2615_;
  assign _1558_ = _0011_[4:2] & _2618_;
  assign _1561_ = _3791_ & _2621_;
  assign _1564_ = _3793_ & _2624_;
  assign _1567_ = { csr_wdata_int_t0[31], csr_wdata_int_t0[4:0] } & _2627_;
  assign _1570_ = csr_mcause_i_t0 & _2630_;
  assign _1575_ = _0035_ & _2635_;
  assign _1580_ = priv_mode_id_o_t0 & _2638_;
  assign _1583_ = mstatus_q_t0[5] & _2633_;
  assign _1588_ = csr_mtval_i_t0 & _2635_;
  assign _1593_ = _0005_ & _2643_;
  assign _1595_ = { csr_wdata_int_t0[31:1], 1'h0 } & _2645_;
  assign _1598_ = _0003_ & _2643_;
  assign _1600_ = _0001_[8:6] & _2648_;
  assign _1603_ = _0001_[1:0] & _2651_;
  assign _1606_ = debug_mode_i_t0 & _2643_;
  assign _1608_ = _0102_ & _2643_;
  assign _1611_ = _0076_ & _2645_;
  assign _1614_ = _0094_ & _2643_;
  assign _1617_ = _0069_ & _2657_;
  assign _1620_ = _0096_ & _2643_;
  assign _1623_ = _0071_ & _2645_;
  assign _1626_ = _0100_ & _2643_;
  assign _1629_ = _0110_ & _2663_;
  assign _1632_ = pc_id_i_t0 & _2666_;
  assign _1635_ = _3795_ & _2669_;
  assign _1638_ = _3797_ & _2672_;
  assign _1643_ = _0005_ & _2607_;
  assign _1646_ = { csr_wdata_int_t0[31:1], 1'h0 } & _2676_;
  assign _1649_ = _0003_ & _2607_;
  assign _1652_ = _0001_[8:6] & _2624_;
  assign _1655_ = _0001_[1:0] & _2681_;
  assign _1658_ = _0015_ & _2607_;
  assign _1661_ = csr_wdata_int_t0 & _2676_;
  assign _1664_ = _0007_ & _2601_;
  assign _1667_ = _3799_ & _2604_;
  assign _1670_ = _3801_ & _2607_;
  assign _1673_ = { csr_wdata_int_t0[31], csr_wdata_int_t0[4:0] } & _2689_;
  assign _1676_ = _3803_ & _2692_;
  assign _1679_ = _3805_ & _2695_;
  assign _1682_ = _0009_ & _2601_;
  assign _1685_ = _3807_ & _2604_;
  assign _1688_ = _3809_ & _2607_;
  assign _1691_ = { csr_wdata_int_t0[31:1], 1'h0 } & _2701_;
  assign _1694_ = _3811_ & _2704_;
  assign _1697_ = _3813_ & _2676_;
  assign _1700_ = _0013_ & _2601_;
  assign _1702_ = _3815_ & _2604_;
  assign _1705_ = _3817_ & _2607_;
  assign _1710_ = priv_mode_id_o_t0 & _2710_;
  assign _1713_ = _3819_ & _2713_;
  assign _1716_ = _3821_ & _2681_;
  assign _1719_ = dcsr_q_t0[31:28] & _2717_;
  assign _1722_ = mstatus_q_t0[5:4] & _2720_;
  assign _1725_ = mstatus_q_t0[3:2] & _2720_;
  assign _1728_ = dcsr_q_t0[15] & _2095_;
  assign _1731_ = dcsr_q_t0[14] & _2095_;
  assign _1733_ = dcsr_q_t0[27:16] & _2725_;
  assign _1736_ = mstatus_q_t0[1:0] & _2720_;
  assign _1739_ = dcsr_q_t0[1:0] & _2729_;
  assign _1742_ = dcsr_q_t0[5] & _2095_;
  assign _1744_ = dcsr_q_t0[4] & _2095_;
  assign _1746_ = dcsr_q_t0[3] & _2095_;
  assign _1748_ = dcsr_q_t0[2] & _2095_;
  assign _1751_ = dcsr_q_t0[13:12] & _2729_;
  assign _1754_ = dcsr_q_t0[11] & _2095_;
  assign _1756_ = csr_wdata_int_t0[1:0] & _2734_;
  assign _1759_ = dcsr_q_t0[9] & _2095_;
  assign _1761_ = csr_wdata_int_t0[12:11] & _2737_;
  assign _1764_ = 32'd0 & _2740_;
  assign _1767_ = 32'd0 & _2743_;
  assign _1770_ = dcsr_q_t0[10] & _2095_;
  assign _1772_ = csr_mtvec_init_i_t0 & _2104_;
  assign _1776_ = 32'd0 & _2748_;
  assign _1791_ = dcsr_q_t0 & _2748_;
  assign _1794_ = csr_mtvec_init_i_t0 & _2746_;
  assign _1809_ = mstatus_q_t0 & _2754_;
  assign _1985_ = { csr_wdata_int_t0[31:8], 8'h00 } & _2757_;
  assign _1988_ = priv_mode_id_o_t0 & _2760_;
  assign _0726_ = _0118_ & _2070_;
  assign _0729_ = csr_wdata_i_t0 & _2073_;
  assign _0732_ = \gen_trigger_regs.selected_tmatch_value_t0 [31] & _2076_;
  assign _0735_ = _0017_[31] & _2079_;
  assign _0738_ = _3244_ & _2082_;
  assign _0743_ = dscratch0_q_t0[31] & _2087_;
  assign _0746_ = _3250_ & _2090_;
  assign _0749_ = _3248_ & _2093_;
  assign _0752_ = dcsr_q_t0[31] & _2096_;
  assign _0755_ = mcause_q_t0[5] & _2099_;
  assign _0758_ = _3258_ & _2102_;
  assign _0761_ = csr_mtvec_o_t0[31] & _2105_;
  assign _0763_ = hart_id_i_t0[31] & _2107_;
  assign _0766_ = _3264_ & _2109_;
  assign _0769_ = _3262_ & _2112_;
  assign _0772_ = _3256_ & _2115_;
  assign _0775_ = \gen_trigger_regs.selected_tmatch_value_t0 [10:8] & _2118_;
  assign _0778_ = _0017_[10:8] & _2121_;
  assign _0781_ = _3272_ & _2124_;
  assign _0784_ = mcountinhibit_t0[10:8] & _2127_;
  assign _0787_ = dscratch0_q_t0[10:8] & _2130_;
  assign _0790_ = _3278_ & _2133_;
  assign _0793_ = _3276_ & _2136_;
  assign _0796_ = dcsr_q_t0[10:8] & _2139_;
  assign _0799_ = csr_mepc_o_t0[10:8] & _2142_;
  assign _0802_ = _3286_ & _2145_;
  assign _0805_ = mscratch_q_t0[10:8] & _2148_;
  assign _0808_ = hart_id_i_t0[10:8] & _2151_;
  assign _0811_ = _3292_ & _2154_;
  assign _0814_ = _3290_ & _2157_;
  assign _0817_ = _3284_ & _2160_;
  assign _0820_ = \gen_trigger_regs.selected_tmatch_value_t0 [7] & _2076_;
  assign _0823_ = _0017_[7] & _2079_;
  assign _0826_ = _3300_ & _2082_;
  assign _0829_ = mcountinhibit_t0[7] & _2085_;
  assign _0832_ = csr_depc_o_t0[7] & _2167_;
  assign _0835_ = dscratch0_q_t0[7] & _2087_;
  assign _0838_ = _3306_ & _2090_;
  assign _0841_ = _3304_ & _2093_;
  assign _0844_ = irq_timer_i_t0 & _2173_;
  assign _0847_ = csr_mepc_o_t0[7] & _2176_;
  assign _0850_ = _3316_ & _2179_;
  assign _0853_ = mscratch_q_t0[7] & _2182_;
  assign _0855_ = hart_id_i_t0[7] & _2107_;
  assign _0858_ = mstatus_q_t0[4] & _2185_;
  assign _0861_ = _3322_ & _2188_;
  assign _0864_ = _3320_ & _2191_;
  assign _0867_ = _3314_ & _2194_;
  assign _0870_ = { 1'h0, cpuctrl_q_t0[5:4] } & _2197_;
  assign _0873_ = 3'h0 & _2200_;
  assign _0876_ = _3332_ & _2203_;
  assign _0879_ = _0017_[6:4] & _2121_;
  assign _0882_ = dscratch1_q_t0[6:4] & _2207_;
  assign _0885_ = mcountinhibit_t0[6:4] & _2127_;
  assign _0888_ = _3338_ & _2211_;
  assign _0891_ = _3336_ & _2214_;
  assign _0894_ = csr_depc_o_t0[6:4] & _2217_;
  assign _0897_ = mtval_q_t0[6:4] & _2220_;
  assign _0900_ = _3348_ & _2223_;
  assign _0903_ = csr_mepc_o_t0[6:4] & _2142_;
  assign _0905_ = hart_id_i_t0[6:4] & _2151_;
  assign _0908_ = mscratch_q_t0[6:4] & _2148_;
  assign _0911_ = _3354_ & _2229_;
  assign _0914_ = _3352_ & _2232_;
  assign _0917_ = _3346_ & _2235_;
  assign _0920_ = 32'd0 & _2238_;
  assign _0923_ = 32'd0 & _2241_;
  assign _0926_ = 32'd0 & _2244_;
  assign _0929_ = 32'd0 & _2247_;
  assign _0932_ = _3365_ & _2250_;
  assign _0935_ = 32'd0 & _2253_;
  assign _0938_ = 32'd0 & _2256_;
  assign _0941_ = 32'd0 & _2259_;
  assign _0944_ = 32'd0 & _2262_;
  assign _0947_ = _3377_ & _2265_;
  assign _0950_ = _3375_ & _2268_;
  assign _0953_ = _3371_ & _2271_;
  assign _0956_ = cpuctrl_q_t0[3] & _2274_;
  assign _0959_ = _0017_[35] & _2277_;
  assign _0964_ = _3385_ & _2281_;
  assign _0967_ = _0019_[3] & _2284_;
  assign _0970_ = dscratch0_q_t0[3] & _2087_;
  assign _0973_ = dscratch1_q_t0[3] & _2288_;
  assign _0976_ = _3393_ & _2291_;
  assign _0979_ = _3391_ & _2294_;
  assign _0982_ = dcsr_q_t0[3] & _2096_;
  assign _0985_ = mcause_q_t0[3] & _2099_;
  assign _0988_ = mtval_q_t0[3] & _2299_;
  assign _0991_ = _3403_ & _2302_;
  assign _0994_ = mscratch_q_t0[3] & _2182_;
  assign _0997_ = csr_mtvec_o_t0[3] & _2105_;
  assign _0999_ = hart_id_i_t0[3] & _2107_;
  assign _1002_ = mstatus_q_t0[5] & _2185_;
  assign _1005_ = _3413_ & _2308_;
  assign _1008_ = _3409_ & _2311_;
  assign _1011_ = _3401_ & _2314_;
  assign _1014_ = \gen_trigger_regs.selected_tmatch_value_t0 [11] & _2076_;
  assign _1017_ = _0017_[11] & _2079_;
  assign _1020_ = _3423_ & _2082_;
  assign _1023_ = mcountinhibit_t0[11] & _2085_;
  assign _1026_ = csr_depc_o_t0[11] & _2167_;
  assign _1029_ = dscratch0_q_t0[11] & _2087_;
  assign _1032_ = _3429_ & _2090_;
  assign _1035_ = _3427_ & _2093_;
  assign _1038_ = irq_external_i_t0 & _2173_;
  assign _1041_ = csr_mepc_o_t0[11] & _2176_;
  assign _1044_ = _3439_ & _2179_;
  assign _1047_ = mscratch_q_t0[11] & _2182_;
  assign _1049_ = hart_id_i_t0[11] & _2107_;
  assign _1052_ = mstatus_q_t0[2] & _2185_;
  assign _1055_ = _3445_ & _2188_;
  assign _1058_ = _3443_ & _2191_;
  assign _1061_ = _3437_ & _2194_;
  assign _1064_ = \gen_trigger_regs.selected_tmatch_value_t0 [21] & _2076_;
  assign _1067_ = _0017_[21] & _2079_;
  assign _1070_ = _3455_ & _2082_;
  assign _1075_ = csr_depc_o_t0[21] & _2167_;
  assign _1078_ = dscratch0_q_t0[21] & _2087_;
  assign _1081_ = _3461_ & _2090_;
  assign _1084_ = _3459_ & _2093_;
  assign _1087_ = irq_fast_i_t0[5] & _2173_;
  assign _1090_ = csr_mepc_o_t0[21] & _2176_;
  assign _1093_ = _3471_ & _2179_;
  assign _1096_ = mscratch_q_t0[21] & _2182_;
  assign _1098_ = hart_id_i_t0[21] & _2107_;
  assign _1101_ = mstatus_q_t0[0] & _2185_;
  assign _1104_ = _3477_ & _2188_;
  assign _1107_ = _3475_ & _2191_;
  assign _1110_ = _3469_ & _2194_;
  assign _1113_ = \mhpmcounter[12]_t0  & _2348_;
  assign _1116_ = 64'h0000000000000000 & _2351_;
  assign _1119_ = \mhpmcounter[9]_t0  & _2354_;
  assign _1122_ = \mhpmcounter[10]_t0  & _2357_;
  assign _1125_ = _3488_ & _2360_;
  assign _1128_ = \mhpmcounter[6]_t0  & _2363_;
  assign _1131_ = \mhpmcounter[7]_t0  & _2366_;
  assign _1134_ = \mhpmcounter[4]_t0  & _2369_;
  assign _1137_ = \mhpmcounter[2]_t0  & _2372_;
  assign _1140_ = _3500_ & _2375_;
  assign _1143_ = _3498_ & _2378_;
  assign _1146_ = _3494_ & _2381_;
  assign _1149_ = \gen_trigger_regs.selected_tmatch_value_t0 [30:22] & _2384_;
  assign _1152_ = _0017_[62:54] & _2387_;
  assign _1155_ = _3508_ & _2390_;
  assign _1158_ = _0019_[30:22] & _2393_;
  assign _1161_ = dscratch0_q_t0[30:22] & _2396_;
  assign _1164_ = dscratch1_q_t0[30:22] & _2399_;
  assign _1167_ = _3514_ & _2402_;
  assign _1170_ = _3512_ & _2405_;
  assign _1173_ = dcsr_q_t0[30:22] & _2408_;
  assign _1176_ = csr_mepc_o_t0[30:22] & _2411_;
  assign _1179_ = mtval_q_t0[30:22] & _2414_;
  assign _1182_ = _3524_ & _2417_;
  assign _1185_ = mscratch_q_t0[30:22] & _2420_;
  assign _1188_ = hart_id_i_t0[30:22] & _2423_;
  assign _1191_ = 9'h000 & _2426_;
  assign _1194_ = _3532_ & _2429_;
  assign _1197_ = _3530_ & _2432_;
  assign _1200_ = _3522_ & _2435_;
  assign _1203_ = _0017_[47:45] & _2438_;
  assign _1206_ = \gen_trigger_regs.selected_tmatch_value_t0 [15:13] & _2118_;
  assign _1209_ = _0019_[15:13] & _2442_;
  assign _1212_ = dscratch1_q_t0[15:13] & _2207_;
  assign _1215_ = _3546_ & _2446_;
  assign _1218_ = _3544_ & _2449_;
  assign _1221_ = csr_depc_o_t0[15:13] & _2217_;
  assign _1224_ = mtval_q_t0[15:13] & _2220_;
  assign _1227_ = _3554_ & _2223_;
  assign _1230_ = csr_mtvec_o_t0[15:13] & _2455_;
  assign _1232_ = hart_id_i_t0[15:13] & _2151_;
  assign _1235_ = _3560_ & _2459_;
  assign _1238_ = _3558_ & _2462_;
  assign _1241_ = _3552_ & _2465_;
  assign _1244_ = \gen_trigger_regs.selected_tmatch_value_t0 [20:18] & _2118_;
  assign _1247_ = _0017_[20:18] & _2121_;
  assign _1250_ = _3568_ & _2124_;
  assign _1253_ = 3'h0 & _2127_;
  assign _1256_ = csr_depc_o_t0[20:18] & _2217_;
  assign _1259_ = dscratch0_q_t0[20:18] & _2130_;
  assign _1262_ = _3574_ & _2133_;
  assign _1265_ = _3572_ & _2136_;
  assign _1268_ = irq_fast_i_t0[4:2] & _2476_;
  assign _1271_ = csr_mepc_o_t0[20:18] & _2142_;
  assign _1274_ = _3584_ & _2480_;
  assign _1277_ = mscratch_q_t0[20:18] & _2148_;
  assign _1279_ = hart_id_i_t0[20:18] & _2151_;
  assign _1285_ = _3590_ & _2488_;
  assign _1288_ = _3588_ & _2491_;
  assign _1291_ = _3582_ & _2494_;
  assign _1294_ = \gen_trigger_regs.selected_tmatch_value_t0 [16] & _2076_;
  assign _1297_ = _0017_[16] & _2079_;
  assign _1300_ = _3600_ & _2082_;
  assign _1305_ = dscratch0_q_t0[16] & _2087_;
  assign _1308_ = _3606_ & _2090_;
  assign _1311_ = _3604_ & _2093_;
  assign _1314_ = dcsr_q_t0[16] & _2096_;
  assign _1317_ = mtval_q_t0[16] & _2299_;
  assign _1320_ = _3614_ & _2302_;
  assign _1323_ = csr_mtvec_o_t0[16] & _2105_;
  assign _1325_ = hart_id_i_t0[16] & _2107_;
  assign _1328_ = mie_q_t0[0] & _2507_;
  assign _1331_ = _3620_ & _2109_;
  assign _1334_ = _3618_ & _2511_;
  assign _1337_ = _3612_ & _2115_;
  assign _1340_ = \gen_trigger_regs.selected_tmatch_value_t0 [17] & _2076_;
  assign _1343_ = _0017_[17] & _2079_;
  assign _1346_ = _3630_ & _2082_;
  assign _1351_ = csr_depc_o_t0[17] & _2167_;
  assign _1354_ = dscratch0_q_t0[17] & _2087_;
  assign _1357_ = _3636_ & _2090_;
  assign _1360_ = _3634_ & _2093_;
  assign _1363_ = irq_fast_i_t0[1] & _2173_;
  assign _1366_ = csr_mepc_o_t0[17] & _2176_;
  assign _1369_ = _3646_ & _2179_;
  assign _1372_ = mscratch_q_t0[17] & _2182_;
  assign _1374_ = hart_id_i_t0[17] & _2107_;
  assign _1377_ = mstatus_q_t0[1] & _2185_;
  assign _1380_ = _3652_ & _2188_;
  assign _1383_ = _3650_ & _2191_;
  assign _1386_ = _3644_ & _2194_;
  assign _1389_ = cpuctrl_q_t0[2:0] & _2197_;
  assign _1392_ = { 2'h0, \gen_trigger_regs.tselect_q_t0  } & _2531_;
  assign _1395_ = { \gen_trigger_regs.selected_tmatch_control_t0 , 2'h0 } & _2200_;
  assign _1398_ = _3662_ & _2203_;
  assign _1401_ = _0017_[2:0] & _2121_;
  assign _1404_ = dscratch1_q_t0[2:0] & _2207_;
  assign _1407_ = { mcountinhibit_t0[2], 1'h0, mcountinhibit_t0[0] } & _2127_;
  assign _1410_ = _3670_ & _2211_;
  assign _1413_ = _3668_ & _2540_;
  assign _1416_ = csr_depc_o_t0[2:0] & _2217_;
  assign _1419_ = mcause_q_t0[2:0] & _2544_;
  assign _1422_ = mtval_q_t0[2:0] & _2220_;
  assign _1425_ = _3680_ & _2223_;
  assign _1428_ = csr_mtvec_o_t0[2:0] & _2455_;
  assign _1430_ = hart_id_i_t0[2:0] & _2151_;
  assign _1282_ = 3'h0 & _2485_;
  assign _1435_ = _3688_ & _2459_;
  assign _1438_ = _3686_ & _2553_;
  assign _1441_ = _3678_ & _2556_;
  assign _1443_ = \gen_trigger_regs.selected_tmatch_value_t0 [12] & _2076_;
  assign _1446_ = _0017_[44] & _2277_;
  assign _1449_ = _3698_ & _2560_;
  assign _1452_ = _0019_[12] & _2284_;
  assign _1455_ = dscratch1_q_t0[12] & _2288_;
  assign _1458_ = _3704_ & _2291_;
  assign _1461_ = _3702_ & _2566_;
  assign _1464_ = csr_depc_o_t0[12] & _2167_;
  assign _1467_ = mtval_q_t0[12] & _2299_;
  assign _1470_ = _3712_ & _2571_;
  assign _1473_ = csr_mtvec_o_t0[12] & _2105_;
  assign _1475_ = hart_id_i_t0[12] & _2107_;
  assign _1478_ = mstatus_q_t0[3] & _2185_;
  assign _1481_ = _3718_ & _2109_;
  assign _1484_ = _3716_ & _2577_;
  assign _1487_ = _3710_ & _2580_;
  assign _1489_ = debug_mode_i_t0 & _2582_;
  assign _1538_ = mstatus_q_t0[4] & _2602_;
  assign _1541_ = _0011_[5] & _2605_;
  assign _1544_ = _0098_[3] & _2608_;
  assign _1549_ = mstack_epc_q_t0 & _2613_;
  assign _1554_ = mstack_q_t0[1:0] & _2616_;
  assign _1556_ = mstack_q_t0[2] & _2611_;
  assign _1559_ = _0114_ & _2619_;
  assign _1562_ = _0011_[4:2] & _2622_;
  assign _1565_ = _0098_[2:0] & _2625_;
  assign _1568_ = mstack_cause_q_t0 & _2628_;
  assign _1571_ = { csr_wdata_int_t0[31], csr_wdata_int_t0[4:0] } & _2631_;
  assign _1573_ = _0007_ & _2634_;
  assign _1576_ = { csr_wdata_int_t0[31:1], 1'h0 } & _2636_;
  assign _1578_ = _0009_ & _2634_;
  assign _1581_ = _0011_[3:2] & _2639_;
  assign _1584_ = _0011_[4] & _2634_;
  assign _1586_ = _0013_ & _2634_;
  assign _1589_ = csr_wdata_int_t0 & _2636_;
  assign _1591_ = _0015_ & _2634_;
  assign _1596_ = _0035_ & _2646_;
  assign _1601_ = debug_cause_i_t0 & _2649_;
  assign _1604_ = priv_mode_id_o_t0 & _2652_;
  assign _1609_ = _0015_ & _2644_;
  assign _1612_ = csr_wdata_int_t0 & _2646_;
  assign _1615_ = _0007_ & _2644_;
  assign _1618_ = { csr_wdata_int_t0[31], csr_wdata_int_t0[4:0] } & _2658_;
  assign _1621_ = _0009_ & _2644_;
  assign _1624_ = { csr_wdata_int_t0[31:1], 1'h0 } & _2646_;
  assign _1627_ = _0013_ & _2644_;
  assign _1630_ = _0011_[5:2] & _2664_;
  assign _1633_ = pc_wb_i_t0 & _2667_;
  assign _1636_ = pc_id_i_t0 & _2670_;
  assign _1639_ = pc_if_i_t0 & _2673_;
  assign _1641_ = _0055_ & _2608_;
  assign _1644_ = _0080_ & _2608_;
  assign _1647_ = _0027_ & _2677_;
  assign _1650_ = _0078_ & _2608_;
  assign _1653_ = _0112_ & _2625_;
  assign _1656_ = _0104_ & _2682_;
  assign _1659_ = _0092_ & _2608_;
  assign _1662_ = _0061_ & _2677_;
  assign _1665_ = _0106_ & _2602_;
  assign _1668_ = _0007_ & _2605_;
  assign _1671_ = _0084_ & _2608_;
  assign _1674_ = _0082_ & _2690_;
  assign _1677_ = { csr_wdata_int_t0[31], csr_wdata_int_t0[4:0] } & _2693_;
  assign _1680_ = _0037_ & _2696_;
  assign _1683_ = _0108_ & _2602_;
  assign _1686_ = _0009_ & _2605_;
  assign _1689_ = _0088_ & _2608_;
  assign _1692_ = _0086_ & _2702_;
  assign _1695_ = { csr_wdata_int_t0[31:1], 1'h0 } & _2705_;
  assign _1698_ = _0043_ & _2677_;
  assign _1703_ = _0013_ & _2605_;
  assign _1706_ = _0090_ & _2608_;
  assign _1708_ = _0011_[5] & _2634_;
  assign _1711_ = mstatus_q_t0[3:2] & _2711_;
  assign _1714_ = dcsr_q_t0[1:0] & _2714_;
  assign _1717_ = 2'h0 & _2682_;
  assign _1720_ = 4'h0 & _2718_;
  assign _1723_ = { csr_wdata_int_t0[3], csr_wdata_int_t0[7] } & _2721_;
  assign _1726_ = _0074_ & _2721_;
  assign _1729_ = csr_wdata_int_t0[15] & _2096_;
  assign _1734_ = 12'h000 & _2726_;
  assign _1737_ = { csr_wdata_int_t0[17], csr_wdata_int_t0[21] } & _2721_;
  assign _1740_ = _0067_ & _2730_;
  assign _1749_ = csr_wdata_int_t0[2] & _2096_;
  assign _1752_ = csr_wdata_int_t0[13:12] & _2730_;
  assign _1757_ = 2'h0 & _2735_;
  assign _1762_ = 2'h0 & _2738_;
  assign _1765_ = _3775_ & _2741_;
  assign _1768_ = _3775_ & _2744_;
  assign _1774_ = _0021_ & _2747_;
  assign _1777_ = _0049_ & _2749_;
  assign _1779_ = _0047_ & _2749_;
  assign _1781_ = _0041_ & _2747_;
  assign _1783_ = _0033_ & _2747_;
  assign _1785_ = _0031_ & _2747_;
  assign _1787_ = _0029_ & _2747_;
  assign _1789_ = _0025_ & _2747_;
  assign _1792_ = { _0023_[31:9], dcsr_q_t0[8:6], _0023_[5:0] } & _2749_;
  assign _1795_ = _0065_ & _2747_;
  assign _1797_ = _0063_ & _2747_;
  assign _1799_ = _0039_ & _2747_;
  assign _1801_ = _0045_ & _2747_;
  assign _1803_ = _0053_ & _2747_;
  assign _1805_ = _0051_ & _2747_;
  assign _1807_ = _0059_ & _2747_;
  assign _1810_ = _0057_ & _2755_;
  assign _1986_ = { boot_addr_i_t0[31:8], 8'h00 } & _2758_;
  assign _1989_ = mstatus_q_t0[3:2] & _2761_;
  assign _1991_ = csr_wdata_int_t0[0] & _2763_;
  assign _2071_ = _0725_ | _0726_;
  assign _2074_ = _0728_ | _0729_;
  assign _2077_ = _0731_ | _0732_;
  assign _2080_ = _0734_ | _0735_;
  assign _2083_ = _0737_ | _0738_;
  assign _2088_ = _0742_ | _0743_;
  assign _2091_ = _0745_ | _0746_;
  assign _2094_ = _0748_ | _0749_;
  assign _2097_ = _0751_ | _0752_;
  assign _2100_ = _0754_ | _0755_;
  assign _2103_ = _0757_ | _0758_;
  assign _2106_ = _0760_ | _0761_;
  assign _2110_ = _0765_ | _0766_;
  assign _2113_ = _0768_ | _0769_;
  assign _2116_ = _0771_ | _0772_;
  assign _2119_ = _0774_ | _0775_;
  assign _2122_ = _0777_ | _0778_;
  assign _2125_ = _0780_ | _0781_;
  assign _2128_ = _0783_ | _0784_;
  assign _2131_ = _0786_ | _0787_;
  assign _2134_ = _0789_ | _0790_;
  assign _2137_ = _0792_ | _0793_;
  assign _2140_ = _0795_ | _0796_;
  assign _2143_ = _0798_ | _0799_;
  assign _2146_ = _0801_ | _0802_;
  assign _2149_ = _0804_ | _0805_;
  assign _2152_ = _0807_ | _0808_;
  assign _2155_ = _0810_ | _0811_;
  assign _2158_ = _0813_ | _0814_;
  assign _2161_ = _0816_ | _0817_;
  assign _2162_ = _0819_ | _0820_;
  assign _2163_ = _0822_ | _0823_;
  assign _2164_ = _0825_ | _0826_;
  assign _2165_ = _0828_ | _0829_;
  assign _2168_ = _0831_ | _0832_;
  assign _2169_ = _0834_ | _0835_;
  assign _2170_ = _0837_ | _0838_;
  assign _2171_ = _0840_ | _0841_;
  assign _2174_ = _0843_ | _0844_;
  assign _2177_ = _0846_ | _0847_;
  assign _2180_ = _0849_ | _0850_;
  assign _2183_ = _0852_ | _0853_;
  assign _2186_ = _0857_ | _0858_;
  assign _2189_ = _0860_ | _0861_;
  assign _2192_ = _0863_ | _0864_;
  assign _2195_ = _0866_ | _0867_;
  assign _2198_ = _0869_ | _0870_;
  assign _2201_ = _0872_ | _0873_;
  assign _2204_ = _0875_ | _0876_;
  assign _2205_ = _0878_ | _0879_;
  assign _2208_ = _0881_ | _0882_;
  assign _2209_ = _0884_ | _0885_;
  assign _2212_ = _0887_ | _0888_;
  assign _2215_ = _0890_ | _0891_;
  assign _2218_ = _0893_ | _0894_;
  assign _2221_ = _0896_ | _0897_;
  assign _2224_ = _0899_ | _0900_;
  assign _2225_ = _0902_ | _0903_;
  assign _2226_ = _0807_ | _0905_;
  assign _2227_ = _0907_ | _0908_;
  assign _2230_ = _0910_ | _0911_;
  assign _2233_ = _0913_ | _0914_;
  assign _2236_ = _0916_ | _0917_;
  assign _2239_ = _0919_ | _0920_;
  assign _2242_ = _0922_ | _0923_;
  assign _2245_ = _0925_ | _0926_;
  assign _2248_ = _0928_ | _0929_;
  assign _2251_ = _0931_ | _0932_;
  assign _2254_ = _0934_ | _0935_;
  assign _2257_ = _0937_ | _0938_;
  assign _2260_ = _0940_ | _0941_;
  assign _2263_ = _0943_ | _0944_;
  assign _2266_ = _0946_ | _0947_;
  assign _2269_ = _0949_ | _0950_;
  assign _2272_ = _0952_ | _0953_;
  assign _2275_ = _0955_ | _0956_;
  assign _2278_ = _0958_ | _0959_;
  assign _2282_ = _0963_ | _0964_;
  assign _2285_ = _0966_ | _0967_;
  assign _2286_ = _0969_ | _0970_;
  assign _2289_ = _0972_ | _0973_;
  assign _2292_ = _0975_ | _0976_;
  assign _2295_ = _0978_ | _0979_;
  assign _2296_ = _0981_ | _0982_;
  assign _2297_ = _0984_ | _0985_;
  assign _2300_ = _0987_ | _0988_;
  assign _2303_ = _0990_ | _0991_;
  assign _2304_ = _0993_ | _0994_;
  assign _2305_ = _0996_ | _0997_;
  assign _2306_ = _1001_ | _1002_;
  assign _2309_ = _1004_ | _1005_;
  assign _2312_ = _1007_ | _1008_;
  assign _2315_ = _1010_ | _1011_;
  assign _2316_ = _1013_ | _1014_;
  assign _2317_ = _1016_ | _1017_;
  assign _2318_ = _1019_ | _1020_;
  assign _2319_ = _1022_ | _1023_;
  assign _2320_ = _1025_ | _1026_;
  assign _2321_ = _1028_ | _1029_;
  assign _2322_ = _1031_ | _1032_;
  assign _2323_ = _1034_ | _1035_;
  assign _2324_ = _1037_ | _1038_;
  assign _2325_ = _1040_ | _1041_;
  assign _2326_ = _1043_ | _1044_;
  assign _2327_ = _1046_ | _1047_;
  assign _2328_ = _1051_ | _1052_;
  assign _2329_ = _1054_ | _1055_;
  assign _2330_ = _1057_ | _1058_;
  assign _2331_ = _1060_ | _1061_;
  assign _2332_ = _1063_ | _1064_;
  assign _2333_ = _1066_ | _1067_;
  assign _2334_ = _1069_ | _1070_;
  assign _2335_ = _1074_ | _1075_;
  assign _2336_ = _1077_ | _1078_;
  assign _2337_ = _1080_ | _1081_;
  assign _2338_ = _1083_ | _1084_;
  assign _2339_ = _1086_ | _1087_;
  assign _2340_ = _1089_ | _1090_;
  assign _2341_ = _1092_ | _1093_;
  assign _2342_ = _1095_ | _1096_;
  assign _2343_ = _1100_ | _1101_;
  assign _2344_ = _1103_ | _1104_;
  assign _2345_ = _1106_ | _1107_;
  assign _2346_ = _1109_ | _1110_;
  assign _2349_ = _1112_ | _1113_;
  assign _2352_ = _1115_ | _1116_;
  assign _2355_ = _1118_ | _1119_;
  assign _2358_ = _1121_ | _1122_;
  assign _2361_ = _1124_ | _1125_;
  assign _2364_ = _1127_ | _1128_;
  assign _2367_ = _1130_ | _1131_;
  assign _2370_ = _1133_ | _1134_;
  assign _2373_ = _1136_ | _1137_;
  assign _2376_ = _1139_ | _1140_;
  assign _2379_ = _1142_ | _1143_;
  assign _2382_ = _1145_ | _1146_;
  assign _2385_ = _1148_ | _1149_;
  assign _2388_ = _1151_ | _1152_;
  assign _2391_ = _1154_ | _1155_;
  assign _2394_ = _1157_ | _1158_;
  assign _2397_ = _1160_ | _1161_;
  assign _2400_ = _1163_ | _1164_;
  assign _2403_ = _1166_ | _1167_;
  assign _2406_ = _1169_ | _1170_;
  assign _2409_ = _1172_ | _1173_;
  assign _2412_ = _1175_ | _1176_;
  assign _2415_ = _1178_ | _1179_;
  assign _2418_ = _1181_ | _1182_;
  assign _2421_ = _1184_ | _1185_;
  assign _2424_ = _1187_ | _1188_;
  assign _2427_ = _1190_ | _1191_;
  assign _2430_ = _1193_ | _1194_;
  assign _2433_ = _1196_ | _1197_;
  assign _2436_ = _1199_ | _1200_;
  assign _2439_ = _1202_ | _1203_;
  assign _2440_ = _1205_ | _1206_;
  assign _2443_ = _1208_ | _1209_;
  assign _2444_ = _1211_ | _1212_;
  assign _2447_ = _1214_ | _1215_;
  assign _2450_ = _1217_ | _1218_;
  assign _2451_ = _1220_ | _1221_;
  assign _2452_ = _1223_ | _1224_;
  assign _2453_ = _1226_ | _1227_;
  assign _2456_ = _1229_ | _1230_;
  assign _2457_ = _0807_ | _1232_;
  assign _2460_ = _1234_ | _1235_;
  assign _2463_ = _1237_ | _1238_;
  assign _2466_ = _1240_ | _1241_;
  assign _2467_ = _1243_ | _1244_;
  assign _2468_ = _1246_ | _1247_;
  assign _2469_ = _1249_ | _1250_;
  assign _2470_ = _1252_ | _1253_;
  assign _2471_ = _1255_ | _1256_;
  assign _2472_ = _1258_ | _1259_;
  assign _2473_ = _1261_ | _1262_;
  assign _2474_ = _1264_ | _1265_;
  assign _2477_ = _1267_ | _1268_;
  assign _2478_ = _1270_ | _1271_;
  assign _2481_ = _1273_ | _1274_;
  assign _2482_ = _1276_ | _1277_;
  assign _2483_ = _0807_ | _1279_;
  assign _2486_ = _1281_ | _1282_;
  assign _2489_ = _1284_ | _1285_;
  assign _2492_ = _1287_ | _1288_;
  assign _2495_ = _1290_ | _1291_;
  assign _2496_ = _1293_ | _1294_;
  assign _2497_ = _1296_ | _1297_;
  assign _2498_ = _1299_ | _1300_;
  assign _2499_ = _1304_ | _1305_;
  assign _2500_ = _1307_ | _1308_;
  assign _2501_ = _1310_ | _1311_;
  assign _2502_ = _1313_ | _1314_;
  assign _2503_ = _1316_ | _1317_;
  assign _2504_ = _1319_ | _1320_;
  assign _2505_ = _1322_ | _1323_;
  assign _2508_ = _1327_ | _1328_;
  assign _2509_ = _1330_ | _1331_;
  assign _2512_ = _1333_ | _1334_;
  assign _2513_ = _1336_ | _1337_;
  assign _2514_ = _1339_ | _1340_;
  assign _2515_ = _1342_ | _1343_;
  assign _2516_ = _1345_ | _1346_;
  assign _2517_ = _1350_ | _1351_;
  assign _2518_ = _1353_ | _1354_;
  assign _2519_ = _1356_ | _1357_;
  assign _2520_ = _1359_ | _1360_;
  assign _2521_ = _1362_ | _1363_;
  assign _2522_ = _1365_ | _1366_;
  assign _2523_ = _1368_ | _1369_;
  assign _2524_ = _1371_ | _1372_;
  assign _2525_ = _1376_ | _1377_;
  assign _2526_ = _1379_ | _1380_;
  assign _2527_ = _1382_ | _1383_;
  assign _2528_ = _1385_ | _1386_;
  assign _2529_ = _1388_ | _1389_;
  assign _2532_ = _1391_ | _1392_;
  assign _2533_ = _1394_ | _1395_;
  assign _2534_ = _1397_ | _1398_;
  assign _2535_ = _1400_ | _1401_;
  assign _2536_ = _1403_ | _1404_;
  assign _2537_ = _1406_ | _1407_;
  assign _2538_ = _1409_ | _1410_;
  assign _2541_ = _1412_ | _1413_;
  assign _2542_ = _1415_ | _1416_;
  assign _2545_ = _1418_ | _1419_;
  assign _2546_ = _1421_ | _1422_;
  assign _2547_ = _1424_ | _1425_;
  assign _2548_ = _1427_ | _1428_;
  assign _2549_ = _0807_ | _1430_;
  assign _2550_ = _1432_ | _1282_;
  assign _2551_ = _1434_ | _1435_;
  assign _2554_ = _1437_ | _1438_;
  assign _2557_ = _1440_ | _1441_;
  assign _2558_ = _1445_ | _1446_;
  assign _2561_ = _1448_ | _1449_;
  assign _2562_ = _1451_ | _1452_;
  assign _2563_ = _1454_ | _1455_;
  assign _2564_ = _1457_ | _1458_;
  assign _2567_ = _1460_ | _1461_;
  assign _2568_ = _1463_ | _1464_;
  assign _2569_ = _1466_ | _1467_;
  assign _2572_ = _1469_ | _1470_;
  assign _2573_ = _1472_ | _1473_;
  assign _2574_ = _1477_ | _1478_;
  assign _2575_ = _1480_ | _1481_;
  assign _2578_ = _1483_ | _1484_;
  assign _2581_ = _1486_ | _1487_;
  assign _2603_ = _1537_ | _1538_;
  assign _2606_ = _1540_ | _1541_;
  assign _2609_ = _1543_ | _1544_;
  assign _2614_ = _1548_ | _1549_;
  assign _2617_ = _1553_ | _1554_;
  assign _2620_ = _1558_ | _1559_;
  assign _2623_ = _1561_ | _1562_;
  assign _2626_ = _1564_ | _1565_;
  assign _2629_ = _1567_ | _1568_;
  assign _2632_ = _1570_ | _1571_;
  assign _2637_ = _1575_ | _1576_;
  assign _2640_ = _1580_ | _1581_;
  assign _2641_ = _1583_ | _1584_;
  assign _2642_ = _1588_ | _1589_;
  assign _2647_ = _1595_ | _1596_;
  assign _2650_ = _1600_ | _1601_;
  assign _2653_ = _1603_ | _1604_;
  assign _2654_ = _1608_ | _1609_;
  assign _2655_ = _1611_ | _1612_;
  assign _2656_ = _1614_ | _1615_;
  assign _2659_ = _1617_ | _1618_;
  assign _2660_ = _1620_ | _1621_;
  assign _2661_ = _1623_ | _1624_;
  assign _2662_ = _1626_ | _1627_;
  assign _2665_ = _1629_ | _1630_;
  assign _2668_ = _1632_ | _1633_;
  assign _2671_ = _1635_ | _1636_;
  assign _2674_ = _1638_ | _1639_;
  assign _2675_ = _1643_ | _1644_;
  assign _2678_ = _1646_ | _1647_;
  assign _2679_ = _1649_ | _1650_;
  assign _2680_ = _1652_ | _1653_;
  assign _2683_ = _1655_ | _1656_;
  assign _2684_ = _1658_ | _1659_;
  assign _2685_ = _1661_ | _1662_;
  assign _2686_ = _1664_ | _1665_;
  assign _2687_ = _1667_ | _1668_;
  assign _2688_ = _1670_ | _1671_;
  assign _2691_ = _1673_ | _1674_;
  assign _2694_ = _1676_ | _1677_;
  assign _2697_ = _1679_ | _1680_;
  assign _2698_ = _1682_ | _1683_;
  assign _2699_ = _1685_ | _1686_;
  assign _2700_ = _1688_ | _1689_;
  assign _2703_ = _1691_ | _1692_;
  assign _2706_ = _1694_ | _1695_;
  assign _2707_ = _1697_ | _1698_;
  assign _2708_ = _1702_ | _1703_;
  assign _2709_ = _1705_ | _1706_;
  assign _2712_ = _1710_ | _1711_;
  assign _2715_ = _1713_ | _1714_;
  assign _2716_ = _1716_ | _1717_;
  assign _2719_ = _1719_ | _1720_;
  assign _2722_ = _1722_ | _1723_;
  assign _2723_ = _1725_ | _1726_;
  assign _2724_ = _1728_ | _1729_;
  assign _2727_ = _1733_ | _1734_;
  assign _2728_ = _1736_ | _1737_;
  assign _2731_ = _1739_ | _1740_;
  assign _2732_ = _1748_ | _1749_;
  assign _2733_ = _1751_ | _1752_;
  assign _2736_ = _1756_ | _1757_;
  assign _2739_ = _1761_ | _1762_;
  assign _2742_ = _1764_ | _1765_;
  assign _2745_ = _1767_ | _1768_;
  assign _2750_ = _1776_ | _1777_;
  assign _2751_ = _1776_ | _1779_;
  assign _2752_ = _1791_ | _1792_;
  assign _2753_ = _1794_ | _1795_;
  assign _2756_ = _1809_ | _1810_;
  assign _2759_ = _1985_ | _1986_;
  assign _2762_ = _1988_ | _1989_;
  assign _2765_ = _3780_ ^ _0117_;
  assign _2766_ = _3241_ ^ csr_wdata_i;
  assign _2767_ = _0016_[63] ^ \gen_trigger_regs.selected_tmatch_value [31];
  assign _2768_ = _0018_[31] ^ _0016_[31];
  assign _2769_ = _3245_ ^ _3243_;
  assign _2770_ = csr_depc_o[31] ^ dscratch0_q[31];
  assign _2771_ = _3251_ ^ _3249_;
  assign _2772_ = _3253_ ^ _3247_;
  assign _2773_ = mtval_q[31] ^ dcsr_q[31];
  assign _2774_ = csr_mepc_o[31] ^ mcause_q[5];
  assign _2775_ = _3259_ ^ _3257_;
  assign _2776_ = mscratch_q[31] ^ csr_mtvec_o[31];
  assign _2777_ = _3265_ ^ _3263_;
  assign _2778_ = _3267_ ^ _3261_;
  assign _2779_ = _3269_ ^ _3255_;
  assign _2780_ = _0016_[42:40] ^ \gen_trigger_regs.selected_tmatch_value [10:8];
  assign _2781_ = _0018_[10:8] ^ _0016_[10:8];
  assign _2782_ = _3273_ ^ _3271_;
  assign _2783_ = dscratch1_q[10:8] ^ mcountinhibit[10:8];
  assign _2784_ = csr_depc_o[10:8] ^ dscratch0_q[10:8];
  assign _2785_ = _3279_ ^ _3277_;
  assign _2786_ = _3281_ ^ _3275_;
  assign _2787_ = mtval_q[10:8] ^ dcsr_q[10:8];
  assign _2788_ = csr_mtvec_o[10:8] ^ csr_mepc_o[10:8];
  assign _2789_ = _3287_ ^ _3285_;
  assign _2790_ = 3'h1 ^ mscratch_q[10:8];
  assign _2791_ = _3293_ ^ _3291_;
  assign _2792_ = _3295_ ^ _3289_;
  assign _2793_ = _3297_ ^ _3283_;
  assign _2794_ = _0016_[39] ^ \gen_trigger_regs.selected_tmatch_value [7];
  assign _2795_ = _0018_[7] ^ _0016_[7];
  assign _2796_ = _3301_ ^ _3299_;
  assign _2797_ = dscratch1_q[7] ^ mcountinhibit[7];
  assign _2798_ = dcsr_q[7] ^ csr_depc_o[7];
  assign _2799_ = _3307_ ^ dscratch0_q[7];
  assign _2800_ = _3309_ ^ _3305_;
  assign _2801_ = _3311_ ^ _3303_;
  assign _2802_ = mtval_q[7] ^ irq_timer_i;
  assign _2803_ = csr_mtvec_o[7] ^ csr_mepc_o[7];
  assign _2804_ = _3317_ ^ _3315_;
  assign _2805_ = mie_q[16] ^ mscratch_q[7];
  assign _2806_ = _3323_ ^ mstatus_q[4];
  assign _2807_ = _3325_ ^ _3321_;
  assign _2808_ = _3327_ ^ _3319_;
  assign _2809_ = _3329_ ^ _3313_;
  assign _2810_ = \gen_trigger_regs.selected_tmatch_value [6:4] ^ { 1'h0, cpuctrl_q[5:4] };
  assign _2811_ = _0016_[38:36] ^ 3'h4;
  assign _2812_ = _3333_ ^ _3331_;
  assign _2813_ = _0018_[6:4] ^ _0016_[6:4];
  assign _2814_ = dscratch0_q[6:4] ^ dscratch1_q[6:4];
  assign _2815_ = _3339_ ^ mcountinhibit[6:4];
  assign _2816_ = _3341_ ^ _3337_;
  assign _2817_ = _3343_ ^ _3335_;
  assign _2818_ = dcsr_q[6:4] ^ csr_depc_o[6:4];
  assign _2819_ = { 2'h0, mcause_q[4] } ^ mtval_q[6:4];
  assign _2820_ = _3349_ ^ _3347_;
  assign _2821_ = csr_mtvec_o[6:4] ^ csr_mepc_o[6:4];
  assign _2822_ = _3355_ ^ mscratch_q[6:4];
  assign _2823_ = _3357_ ^ _3353_;
  assign _2824_ = _3359_ ^ _3351_;
  assign _2825_ = _3361_ ^ _3345_;
  assign _2827_ = _3366_ ^ 32'd1024;
  assign _2828_ = _3368_ ^ _3364_;
  assign _2829_ = _3372_ ^ 32'd128;
  assign _2830_ = _3378_ ^ _3376_;
  assign _2831_ = _3380_ ^ _3374_;
  assign _2832_ = _3382_ ^ _3370_;
  assign _2833_ = \gen_trigger_regs.selected_tmatch_value [3] ^ cpuctrl_q[3];
  assign _2834_ = _0016_[3] ^ _0016_[35];
  assign _2835_ = _3388_ ^ _3384_;
  assign _2836_ = mcountinhibit[3] ^ _0018_[3];
  assign _2837_ = csr_depc_o[3] ^ dscratch0_q[3];
  assign _2838_ = _3394_ ^ dscratch1_q[3];
  assign _2839_ = _3396_ ^ _3392_;
  assign _2840_ = _3398_ ^ _3390_;
  assign _2841_ = irq_software_i ^ dcsr_q[3];
  assign _2842_ = csr_mepc_o[3] ^ mcause_q[3];
  assign _2843_ = _3404_ ^ mtval_q[3];
  assign _2844_ = _3406_ ^ _3402_;
  assign _2845_ = mie_q[17] ^ mscratch_q[3];
  assign _2846_ = _3410_ ^ csr_mtvec_o[3];
  assign _2847_ = _3414_ ^ mstatus_q[5];
  assign _2848_ = _3416_ ^ _3412_;
  assign _2849_ = _3418_ ^ _3408_;
  assign _2850_ = _3420_ ^ _3400_;
  assign _2851_ = _0016_[43] ^ \gen_trigger_regs.selected_tmatch_value [11];
  assign _2852_ = _0018_[11] ^ _0016_[11];
  assign _2853_ = _3424_ ^ _3422_;
  assign _2854_ = dscratch1_q[11] ^ mcountinhibit[11];
  assign _2855_ = dcsr_q[11] ^ csr_depc_o[11];
  assign _2856_ = _3430_ ^ dscratch0_q[11];
  assign _2857_ = _3432_ ^ _3428_;
  assign _2858_ = _3434_ ^ _3426_;
  assign _2859_ = mtval_q[11] ^ irq_external_i;
  assign _2860_ = csr_mtvec_o[11] ^ csr_mepc_o[11];
  assign _2861_ = _3440_ ^ _3438_;
  assign _2862_ = mie_q[15] ^ mscratch_q[11];
  assign _2863_ = _3446_ ^ mstatus_q[2];
  assign _2864_ = _3448_ ^ _3444_;
  assign _2865_ = _3450_ ^ _3442_;
  assign _2866_ = _3452_ ^ _3436_;
  assign _2867_ = _0016_[53] ^ \gen_trigger_regs.selected_tmatch_value [21];
  assign _2868_ = _0018_[21] ^ _0016_[21];
  assign _2869_ = _3456_ ^ _3454_;
  assign _2870_ = dcsr_q[21] ^ csr_depc_o[21];
  assign _2871_ = _3462_ ^ dscratch0_q[21];
  assign _2872_ = _3464_ ^ _3460_;
  assign _2873_ = _3466_ ^ _3458_;
  assign _2874_ = mtval_q[21] ^ irq_fast_i[5];
  assign _2875_ = csr_mtvec_o[21] ^ csr_mepc_o[21];
  assign _2876_ = _3472_ ^ _3470_;
  assign _2877_ = mie_q[5] ^ mscratch_q[21];
  assign _2878_ = _3478_ ^ mstatus_q[0];
  assign _2879_ = _3480_ ^ _3476_;
  assign _2880_ = _3482_ ^ _3474_;
  assign _2881_ = _3484_ ^ _3468_;
  assign _2882_ = \mhpmcounter[11]  ^ \mhpmcounter[12] ;
  assign _2884_ = \mhpmcounter[8]  ^ \mhpmcounter[9] ;
  assign _2885_ = _3489_ ^ \mhpmcounter[10] ;
  assign _2886_ = _3491_ ^ _3487_;
  assign _2887_ = \mhpmcounter[5]  ^ \mhpmcounter[6] ;
  assign _2888_ = _3495_ ^ \mhpmcounter[7] ;
  assign _2889_ = \mhpmcounter[3]  ^ \mhpmcounter[4] ;
  assign _2890_ = \mhpmcounter[0]  ^ \mhpmcounter[2] ;
  assign _2891_ = _3501_ ^ _3499_;
  assign _2892_ = _3503_ ^ _3497_;
  assign _2893_ = _3505_ ^ _3493_;
  assign _2894_ = 9'h0a0 ^ \gen_trigger_regs.selected_tmatch_value [30:22];
  assign _2895_ = _0016_[30:22] ^ _0016_[62:54];
  assign _2896_ = _3509_ ^ _3507_;
  assign _2897_ = 9'h1ff ^ _0018_[30:22];
  assign _2898_ = csr_depc_o[30:22] ^ dscratch0_q[30:22];
  assign _2899_ = _3515_ ^ dscratch1_q[30:22];
  assign _2900_ = _3517_ ^ _3513_;
  assign _2901_ = _3519_ ^ _3511_;
  assign _2902_ = irq_fast_i[14:6] ^ dcsr_q[30:22];
  assign _2903_ = csr_mtvec_o[30:22] ^ csr_mepc_o[30:22];
  assign _2904_ = _3525_ ^ mtval_q[30:22];
  assign _2905_ = _3527_ ^ _3523_;
  assign _2906_ = mie_q[14:6] ^ mscratch_q[30:22];
  assign _2907_ = _3533_ ^ 9'h100;
  assign _2908_ = _3535_ ^ _3531_;
  assign _2909_ = _3537_ ^ _3529_;
  assign _2910_ = _3539_ ^ _3521_;
  assign _2911_ = _0016_[15:13] ^ _0016_[47:45];
  assign _2912_ = _3541_ ^ \gen_trigger_regs.selected_tmatch_value [15:13];
  assign _2913_ = 3'h7 ^ _0018_[15:13];
  assign _2914_ = dscratch0_q[15:13] ^ dscratch1_q[15:13];
  assign _2915_ = _3547_ ^ _3545_;
  assign _2916_ = _3549_ ^ _3543_;
  assign _2917_ = dcsr_q[15:13] ^ csr_depc_o[15:13];
  assign _2918_ = csr_mepc_o[15:13] ^ mtval_q[15:13];
  assign _2919_ = _3555_ ^ _3553_;
  assign _2920_ = mscratch_q[15:13] ^ csr_mtvec_o[15:13];
  assign _2921_ = _3561_ ^ _3559_;
  assign _2922_ = _3563_ ^ _3557_;
  assign _2923_ = _3565_ ^ _3551_;
  assign _2924_ = _0016_[52:50] ^ \gen_trigger_regs.selected_tmatch_value [20:18];
  assign _2925_ = _0018_[20:18] ^ _0016_[20:18];
  assign _2926_ = _3569_ ^ _3567_;
  assign _2927_ = dscratch1_q[20:18] ^ 3'h7;
  assign _2928_ = dcsr_q[20:18] ^ csr_depc_o[20:18];
  assign _2929_ = _3575_ ^ dscratch0_q[20:18];
  assign _2930_ = _3577_ ^ _3573_;
  assign _2931_ = _3579_ ^ _3571_;
  assign _2932_ = mtval_q[20:18] ^ irq_fast_i[4:2];
  assign _2933_ = csr_mtvec_o[20:18] ^ csr_mepc_o[20:18];
  assign _2934_ = _3585_ ^ _3583_;
  assign _2935_ = mie_q[4:2] ^ mscratch_q[20:18];
  assign _2936_ = _3591_ ^ 3'h4;
  assign _2937_ = _3593_ ^ _3589_;
  assign _2938_ = _3595_ ^ _3587_;
  assign _2939_ = _3597_ ^ _3581_;
  assign _2940_ = _0016_[48] ^ \gen_trigger_regs.selected_tmatch_value [16];
  assign _2941_ = _0018_[16] ^ _0016_[16];
  assign _2942_ = _3601_ ^ _3599_;
  assign _2943_ = csr_depc_o[16] ^ dscratch0_q[16];
  assign _2944_ = _3607_ ^ _3605_;
  assign _2945_ = _3609_ ^ _3603_;
  assign _2946_ = irq_fast_i[0] ^ dcsr_q[16];
  assign _2947_ = csr_mepc_o[16] ^ mtval_q[16];
  assign _2948_ = _3615_ ^ _3613_;
  assign _2949_ = mscratch_q[16] ^ csr_mtvec_o[16];
  assign _2950_ = _3621_ ^ mie_q[0];
  assign _2951_ = _3623_ ^ _3619_;
  assign _2952_ = _3625_ ^ _3617_;
  assign _2953_ = _3627_ ^ _3611_;
  assign _2954_ = _0016_[49] ^ \gen_trigger_regs.selected_tmatch_value [17];
  assign _2955_ = _0018_[17] ^ _0016_[17];
  assign _2956_ = _3631_ ^ _3629_;
  assign _2957_ = dcsr_q[17] ^ csr_depc_o[17];
  assign _2958_ = _3637_ ^ dscratch0_q[17];
  assign _2959_ = _3639_ ^ _3635_;
  assign _2960_ = _3641_ ^ _3633_;
  assign _2961_ = mtval_q[17] ^ irq_fast_i[1];
  assign _2962_ = csr_mtvec_o[17] ^ csr_mepc_o[17];
  assign _2963_ = _3647_ ^ _3645_;
  assign _2964_ = mie_q[1] ^ mscratch_q[17];
  assign _2965_ = _3653_ ^ mstatus_q[1];
  assign _2966_ = _3655_ ^ _3651_;
  assign _2967_ = _3657_ ^ _3649_;
  assign _2968_ = _3659_ ^ _3643_;
  assign _2969_ = \gen_trigger_regs.selected_tmatch_value [2:0] ^ cpuctrl_q[2:0];
  assign _2970_ = _0016_[34:32] ^ { 2'h0, \gen_trigger_regs.tselect_q  };
  assign _2971_ = _3663_ ^ { \gen_trigger_regs.selected_tmatch_control , 2'h0 };
  assign _2972_ = _3665_ ^ _3661_;
  assign _2973_ = _0018_[2:0] ^ _0016_[2:0];
  assign _2974_ = dscratch0_q[2:0] ^ dscratch1_q[2:0];
  assign _2975_ = _3671_ ^ { mcountinhibit[2], 1'h0, mcountinhibit[0] };
  assign _2976_ = _3673_ ^ _3669_;
  assign _2977_ = _3675_ ^ _3667_;
  assign _2978_ = dcsr_q[2:0] ^ csr_depc_o[2:0];
  assign _2979_ = csr_mepc_o[2:0] ^ mcause_q[2:0];
  assign _2980_ = _3681_ ^ mtval_q[2:0];
  assign _2981_ = _3683_ ^ _3679_;
  assign _2982_ = mscratch_q[2:0] ^ csr_mtvec_o[2:0];
  assign _2983_ = _3689_ ^ 3'h4;
  assign _2984_ = _3691_ ^ _3687_;
  assign _2985_ = _3693_ ^ _3685_;
  assign _2986_ = _3695_ ^ _3677_;
  assign _2987_ = _0016_[12] ^ _0016_[44];
  assign _2988_ = _3699_ ^ _3697_;
  assign _2989_ = mcountinhibit[12] ^ _0018_[12];
  assign _2990_ = dscratch0_q[12] ^ dscratch1_q[12];
  assign _2991_ = _3705_ ^ _3703_;
  assign _2992_ = _3707_ ^ _3701_;
  assign _2993_ = dcsr_q[12] ^ csr_depc_o[12];
  assign _2994_ = csr_mepc_o[12] ^ mtval_q[12];
  assign _2995_ = _3713_ ^ _3711_;
  assign _2996_ = mscratch_q[12] ^ csr_mtvec_o[12];
  assign _2997_ = _3719_ ^ mstatus_q[3];
  assign _2998_ = _3721_ ^ _3717_;
  assign _2999_ = _3723_ ^ _3715_;
  assign _3000_ = _3725_ ^ _3709_;
  assign _3003_ = _0010_[5] ^ mstatus_q[4];
  assign _3004_ = _3786_ ^ _0010_[5];
  assign _3005_ = _3788_ ^ _0097_[3];
  assign _3006_ = { csr_wdata_int[31:1], 1'h0 } ^ mstack_epc_q;
  assign _3007_ = _0010_[4:2] ^ _0113_;
  assign _3008_ = _3790_ ^ _0010_[4:2];
  assign _3009_ = _3792_ ^ _0097_[2:0];
  assign _3010_ = { csr_wdata_int[31], csr_wdata_int[4:0] } ^ mstack_cause_q;
  assign _3011_ = csr_mcause_i ^ { csr_wdata_int[31], csr_wdata_int[4:0] };
  assign _3013_ = priv_mode_id_o ^ _0010_[3:2];
  assign _3014_ = mstatus_q[5] ^ _0010_[4];
  assign _3015_ = csr_mtval_i ^ csr_wdata_int;
  assign _3012_ = { csr_wdata_int[31:1], 1'h0 } ^ _0034_;
  assign _3016_ = _0000_[8:6] ^ debug_cause_i;
  assign _3017_ = _0000_[1:0] ^ priv_mode_id_o;
  assign _3018_ = _0101_ ^ _0014_;
  assign _3019_ = _0075_ ^ csr_wdata_int;
  assign _3020_ = _0093_ ^ _0006_;
  assign _3021_ = _0068_ ^ { csr_wdata_int[31], csr_wdata_int[4:0] };
  assign _3022_ = _0095_ ^ _0008_;
  assign _3023_ = _0070_ ^ { csr_wdata_int[31:1], 1'h0 };
  assign _3024_ = _0099_ ^ _0012_;
  assign _3025_ = _0109_ ^ _0010_[5:2];
  assign _3026_ = pc_id_i ^ pc_wb_i;
  assign _3027_ = _3794_ ^ pc_id_i;
  assign _3028_ = _3796_ ^ pc_if_i;
  assign _3029_ = _0004_ ^ _0079_;
  assign _3030_ = { csr_wdata_int[31:1], 1'h0 } ^ _0026_;
  assign _3031_ = _0002_ ^ _0077_;
  assign _3032_ = _0000_[8:6] ^ _0111_;
  assign _3033_ = _0000_[1:0] ^ _0103_;
  assign _3034_ = _0014_ ^ _0091_;
  assign _3035_ = csr_wdata_int ^ _0060_;
  assign _3036_ = _0006_ ^ _0105_;
  assign _3037_ = _3798_ ^ _0006_;
  assign _3038_ = _3800_ ^ _0083_;
  assign _3039_ = { csr_wdata_int[31], csr_wdata_int[4:0] } ^ _0081_;
  assign _3040_ = _3802_ ^ { csr_wdata_int[31], csr_wdata_int[4:0] };
  assign _3041_ = _3804_ ^ _0036_;
  assign _3042_ = _0008_ ^ _0107_;
  assign _3043_ = _3806_ ^ _0008_;
  assign _3044_ = _3808_ ^ _0087_;
  assign _3045_ = { csr_wdata_int[31:1], 1'h0 } ^ _0085_;
  assign _3046_ = _3810_ ^ { csr_wdata_int[31:1], 1'h0 };
  assign _3047_ = _3812_ ^ _0042_;
  assign _3048_ = _3814_ ^ _0012_;
  assign _3049_ = _3816_ ^ _0089_;
  assign _3050_ = priv_mode_id_o ^ mstatus_q[3:2];
  assign _3051_ = _3818_ ^ dcsr_q[1:0];
  assign _3052_ = _3820_ ^ 2'h3;
  assign _3053_ = dcsr_q[31:28] ^ 4'h4;
  assign _3054_ = mstatus_q[5:4] ^ { csr_wdata_int[3], csr_wdata_int[7] };
  assign _3055_ = mstatus_q[3:2] ^ _0073_;
  assign _3056_ = dcsr_q[15] ^ csr_wdata_int[15];
  assign _3057_ = mstatus_q[1:0] ^ { csr_wdata_int[17], csr_wdata_int[21] };
  assign _3058_ = dcsr_q[1:0] ^ _0066_;
  assign _3059_ = dcsr_q[2] ^ csr_wdata_int[2];
  assign _3060_ = dcsr_q[13:12] ^ csr_wdata_int[13:12];
  assign _3061_ = csr_wdata_int[1:0] ^ 2'h3;
  assign _3062_ = csr_wdata_int[12:11] ^ 2'h3;
  assign _3064_ = dcsr_q ^ { _0022_[31:9], dcsr_q[8:6], _0022_[5:0] };
  assign _3065_ = csr_mtvec_init_i ^ _0064_;
  assign _3066_ = mstatus_q ^ _0056_;
  assign _3067_ = { csr_wdata_int[31:8], 8'h01 } ^ { boot_addr_i[31:8], 8'h01 };
  assign _0727_ = { _3732_, _3732_, _3732_, _3732_, _3732_, _3732_, _3732_, _3732_, _3732_, _3732_, _3732_, _3732_, _3732_, _3732_, _3732_, _3732_, _3732_, _3732_, _3732_, _3732_, _3732_, _3732_, _3732_, _3732_, _3732_, _3732_, _3732_, _3732_, _3732_, _3732_, _3732_, _3732_ } & _2765_;
  assign _0730_ = { _0161_, _0161_, _0161_, _0161_, _0161_, _0161_, _0161_, _0161_, _0161_, _0161_, _0161_, _0161_, _0161_, _0161_, _0161_, _0161_, _0161_, _0161_, _0161_, _0161_, _0161_, _0161_, _0161_, _0161_, _0161_, _0161_, _0161_, _0161_, _0161_, _0161_, _0161_, _0161_ } & _2766_;
  assign _0733_ = _3743_ & _2767_;
  assign _0736_ = _3831_ & _2768_;
  assign _0739_ = _1994_ & _2769_;
  assign _0741_ = _0041_ & _0412_;
  assign _0744_ = _0031_ & _2770_;
  assign _0747_ = _1996_ & _2771_;
  assign _0750_ = _0429_ & _2772_;
  assign _0753_ = _0025_ & _2773_;
  assign _0756_ = _0039_ & _2774_;
  assign _0759_ = _1998_ & _2775_;
  assign _0762_ = _3838_ & _2776_;
  assign _0764_ = _3889_ & hart_id_i[31];
  assign _0767_ = _2000_ & _2777_;
  assign _0770_ = _0431_ & _2778_;
  assign _0773_ = _0433_ & _2779_;
  assign _0776_ = { _3743_, _3743_, _3743_ } & _2780_;
  assign _0779_ = { _3831_, _3831_, _3831_ } & _2781_;
  assign _0782_ = { _1994_, _1994_, _1994_ } & _2782_;
  assign _0785_ = { _0041_, _0041_, _0041_ } & _2783_;
  assign _0788_ = { _0031_, _0031_, _0031_ } & _2784_;
  assign _0791_ = { _1996_, _1996_, _1996_ } & _2785_;
  assign _0794_ = { _0429_, _0429_, _0429_ } & _2786_;
  assign _0797_ = { _0025_, _0025_, _0025_ } & _2787_;
  assign _0800_ = { _0045_, _0045_, _0045_ } & _2788_;
  assign _0803_ = { _1998_, _1998_, _1998_ } & _2789_;
  assign _0806_ = { _0053_, _0053_, _0053_ } & _2790_;
  assign _0809_ = { _3889_, _3889_, _3889_ } & hart_id_i[10:8];
  assign _0812_ = { _2002_, _2002_, _2002_ } & _2791_;
  assign _0815_ = { _0435_, _0435_, _0435_ } & _2792_;
  assign _0818_ = { _0433_, _0433_, _0433_ } & _2793_;
  assign _0821_ = _3743_ & _2794_;
  assign _0824_ = _3831_ & _2795_;
  assign _0827_ = _1994_ & _2796_;
  assign _0830_ = _0041_ & _2797_;
  assign _0833_ = _0029_ & _2798_;
  assign _0836_ = _0031_ & _2799_;
  assign _0839_ = _1996_ & _2800_;
  assign _0842_ = _0429_ & _2801_;
  assign _0845_ = _3893_ & _2802_;
  assign _0848_ = _0045_ & _2803_;
  assign _0851_ = _2004_ & _2804_;
  assign _0854_ = _0053_ & _2805_;
  assign _0856_ = _3889_ & hart_id_i[7];
  assign _0859_ = _0059_ & _2806_;
  assign _0862_ = _2006_ & _2807_;
  assign _0865_ = _0437_ & _2808_;
  assign _0868_ = _0439_ & _2809_;
  assign _0871_ = { _0021_, _0021_, _0021_ } & _2810_;
  assign _0874_ = { _3741_, _3741_, _3741_ } & _2811_;
  assign _0877_ = { _2008_, _2008_, _2008_ } & _2812_;
  assign _0880_ = { _3831_, _3831_, _3831_ } & _2813_;
  assign _0883_ = { _0033_, _0033_, _0033_ } & _2814_;
  assign _0886_ = { _0041_, _0041_, _0041_ } & _2815_;
  assign _0889_ = { _2010_, _2010_, _2010_ } & _2816_;
  assign _0892_ = { _0441_, _0441_, _0441_ } & _2817_;
  assign _0895_ = { _0029_, _0029_, _0029_ } & _2818_;
  assign _0898_ = { _0063_, _0063_, _0063_ } & _2819_;
  assign _0901_ = { _2012_, _2012_, _2012_ } & _2820_;
  assign _0904_ = { _0045_, _0045_, _0045_ } & _2821_;
  assign _0906_ = { _3889_, _3889_, _3889_ } & hart_id_i[6:4];
  assign _0909_ = { _0053_, _0053_, _0053_ } & _2822_;
  assign _0912_ = { _2014_, _2014_, _2014_ } & _2823_;
  assign _0915_ = { _0443_, _0443_, _0443_ } & _2824_;
  assign _0918_ = { _0445_, _0445_, _0445_ } & _2825_;
  assign _0921_ = { _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_ } & 32'd6144;
  assign _0924_ = { _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_ } & _2826_;
  assign _0927_ = { _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_ } & 32'd768;
  assign _0930_ = { _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_ } & _2827_;
  assign _0933_ = { _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_ } & _2828_;
  assign _0936_ = { _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_ } & 32'd96;
  assign _0939_ = { _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_ } & _2829_;
  assign _0942_ = { _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_ } & 32'd24;
  assign _0945_ = { _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_ } & 32'd5;
  assign _0948_ = { _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_ } & _2830_;
  assign _0951_ = { _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_ } & _2831_;
  assign _0954_ = { _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_ } & _2832_;
  assign _0957_ = _0021_ & _2833_;
  assign _0960_ = _3827_ & _2834_;
  assign _0962_ = _3741_ & _0413_;
  assign _0965_ = _2008_ & _2835_;
  assign _0968_ = _3847_ & _2836_;
  assign _0971_ = _0031_ & _2837_;
  assign _0974_ = _0033_ & _2838_;
  assign _0977_ = _2018_ & _2839_;
  assign _0980_ = _0453_ & _2840_;
  assign _0983_ = _0025_ & _2841_;
  assign _0986_ = _0039_ & _2842_;
  assign _0989_ = _0063_ & _2843_;
  assign _0992_ = _2020_ & _2844_;
  assign _0995_ = _0053_ & _2845_;
  assign _0998_ = _3838_ & _2846_;
  assign _1000_ = _3889_ & hart_id_i[3];
  assign _1003_ = _0059_ & _2847_;
  assign _1006_ = _0455_ & _2848_;
  assign _1009_ = _0457_ & _2849_;
  assign _1012_ = _0459_ & _2850_;
  assign _1015_ = _3743_ & _2851_;
  assign _1018_ = _3831_ & _2852_;
  assign _1021_ = _1994_ & _2853_;
  assign _1024_ = _0041_ & _2854_;
  assign _1027_ = _0029_ & _2855_;
  assign _1030_ = _0031_ & _2856_;
  assign _1033_ = _1996_ & _2857_;
  assign _1036_ = _0429_ & _2858_;
  assign _1039_ = _3893_ & _2859_;
  assign _1042_ = _0045_ & _2860_;
  assign _1045_ = _2004_ & _2861_;
  assign _1048_ = _0053_ & _2862_;
  assign _1050_ = _3889_ & hart_id_i[11];
  assign _1053_ = _0059_ & _2863_;
  assign _1056_ = _2006_ & _2864_;
  assign _1059_ = _0437_ & _2865_;
  assign _1062_ = _0439_ & _2866_;
  assign _1065_ = _3743_ & _2867_;
  assign _1068_ = _3831_ & _2868_;
  assign _1071_ = _1994_ & _2869_;
  assign _1073_ = _0041_ & _0414_;
  assign _1076_ = _0029_ & _2870_;
  assign _1079_ = _0031_ & _2871_;
  assign _1082_ = _1996_ & _2872_;
  assign _1085_ = _0429_ & _2873_;
  assign _1088_ = _3893_ & _2874_;
  assign _1091_ = _0045_ & _2875_;
  assign _1094_ = _2004_ & _2876_;
  assign _1097_ = _0053_ & _2877_;
  assign _1099_ = _3889_ & hart_id_i[21];
  assign _1102_ = _0059_ & _2878_;
  assign _1105_ = _2006_ & _2879_;
  assign _1108_ = _0437_ & _2880_;
  assign _1111_ = _0439_ & _2881_;
  assign _1114_ = { _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_, _3933_ } & _2882_;
  assign _1117_ = { _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_, _0155_ } & _2883_;
  assign _1120_ = { _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_, _3939_ } & _2884_;
  assign _1123_ = { _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_, _3937_ } & _2885_;
  assign _1126_ = { _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_ } & _2886_;
  assign _1129_ = { _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_, _3945_ } & _2887_;
  assign _1132_ = { _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_, _3943_ } & _2888_;
  assign _1135_ = { _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_, _3949_ } & _2889_;
  assign _1138_ = { _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_, _3953_ } & _2890_;
  assign _1141_ = { _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_, _2016_ } & _2891_;
  assign _1144_ = { _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_ } & _2892_;
  assign _1147_ = { _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_, _0451_ } & _2893_;
  assign _1150_ = { _3743_, _3743_, _3743_, _3743_, _3743_, _3743_, _3743_, _3743_, _3743_ } & _2894_;
  assign _1153_ = { _3827_, _3827_, _3827_, _3827_, _3827_, _3827_, _3827_, _3827_, _3827_ } & _2895_;
  assign _1156_ = { _2022_, _2022_, _2022_, _2022_, _2022_, _2022_, _2022_, _2022_, _2022_ } & _2896_;
  assign _1159_ = { _3847_, _3847_, _3847_, _3847_, _3847_, _3847_, _3847_, _3847_, _3847_ } & _2897_;
  assign _1162_ = { _0031_, _0031_, _0031_, _0031_, _0031_, _0031_, _0031_, _0031_, _0031_ } & _2898_;
  assign _1165_ = { _0033_, _0033_, _0033_, _0033_, _0033_, _0033_, _0033_, _0033_, _0033_ } & _2899_;
  assign _1168_ = { _2018_, _2018_, _2018_, _2018_, _2018_, _2018_, _2018_, _2018_, _2018_ } & _2900_;
  assign _1171_ = { _0461_, _0461_, _0461_, _0461_, _0461_, _0461_, _0461_, _0461_, _0461_ } & _2901_;
  assign _1174_ = { _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_ } & _2902_;
  assign _1177_ = { _0045_, _0045_, _0045_, _0045_, _0045_, _0045_, _0045_, _0045_, _0045_ } & _2903_;
  assign _1180_ = { _0063_, _0063_, _0063_, _0063_, _0063_, _0063_, _0063_, _0063_, _0063_ } & _2904_;
  assign _1183_ = { _2020_, _2020_, _2020_, _2020_, _2020_, _2020_, _2020_, _2020_, _2020_ } & _2905_;
  assign _1186_ = { _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_ } & _2906_;
  assign _1189_ = { _3889_, _3889_, _3889_, _3889_, _3889_, _3889_, _3889_, _3889_, _3889_ } & hart_id_i[30:22];
  assign _1192_ = { _3891_, _3891_, _3891_, _3891_, _3891_, _3891_, _3891_, _3891_, _3891_ } & _2907_;
  assign _1195_ = { _2006_, _2006_, _2006_, _2006_, _2006_, _2006_, _2006_, _2006_, _2006_ } & _2908_;
  assign _1198_ = { _0463_, _0463_, _0463_, _0463_, _0463_, _0463_, _0463_, _0463_, _0463_ } & _2909_;
  assign _1201_ = { _0465_, _0465_, _0465_, _0465_, _0465_, _0465_, _0465_, _0465_, _0465_ } & _2910_;
  assign _1204_ = { _3827_, _3827_, _3827_ } & _2911_;
  assign _1207_ = { _3743_, _3743_, _3743_ } & _2912_;
  assign _1210_ = { _3847_, _3847_, _3847_ } & _2913_;
  assign _1213_ = { _0033_, _0033_, _0033_ } & _2914_;
  assign _1216_ = { _2018_, _2018_, _2018_ } & _2915_;
  assign _1219_ = { _0467_, _0467_, _0467_ } & _2916_;
  assign _1222_ = { _0029_, _0029_, _0029_ } & _2917_;
  assign _1225_ = { _0063_, _0063_, _0063_ } & _2918_;
  assign _1228_ = { _2012_, _2012_, _2012_ } & _2919_;
  assign _1231_ = { _3838_, _3838_, _3838_ } & _2920_;
  assign _1233_ = { _3889_, _3889_, _3889_ } & hart_id_i[15:13];
  assign _1236_ = { _2000_, _2000_, _2000_ } & _2921_;
  assign _1239_ = { _0469_, _0469_, _0469_ } & _2922_;
  assign _1242_ = { _0471_, _0471_, _0471_ } & _2923_;
  assign _1245_ = { _3743_, _3743_, _3743_ } & _2924_;
  assign _1248_ = { _3831_, _3831_, _3831_ } & _2925_;
  assign _1251_ = { _1994_, _1994_, _1994_ } & _2926_;
  assign _1254_ = { _0041_, _0041_, _0041_ } & _2927_;
  assign _1257_ = { _0029_, _0029_, _0029_ } & _2928_;
  assign _1260_ = { _0031_, _0031_, _0031_ } & _2929_;
  assign _1263_ = { _1996_, _1996_, _1996_ } & _2930_;
  assign _1266_ = { _0429_, _0429_, _0429_ } & _2931_;
  assign _1269_ = { _3893_, _3893_, _3893_ } & _2932_;
  assign _1272_ = { _0045_, _0045_, _0045_ } & _2933_;
  assign _1275_ = { _2004_, _2004_, _2004_ } & _2934_;
  assign _1278_ = { _0053_, _0053_, _0053_ } & _2935_;
  assign _1280_ = { _3889_, _3889_, _3889_ } & hart_id_i[20:18];
  assign _1283_ = { _3891_, _3891_, _3891_ } & _2936_;
  assign _1286_ = { _2006_, _2006_, _2006_ } & _2937_;
  assign _1289_ = { _0437_, _0437_, _0437_ } & _2938_;
  assign _1292_ = { _0439_, _0439_, _0439_ } & _2939_;
  assign _1295_ = _3743_ & _2940_;
  assign _1298_ = _3831_ & _2941_;
  assign _1301_ = _1994_ & _2942_;
  assign _1303_ = _0041_ & _0415_;
  assign _1306_ = _0031_ & _2943_;
  assign _1309_ = _1996_ & _2944_;
  assign _1312_ = _0429_ & _2945_;
  assign _1315_ = _0025_ & _2946_;
  assign _1318_ = _0063_ & _2947_;
  assign _1321_ = _2020_ & _2948_;
  assign _1324_ = _3838_ & _2949_;
  assign _1326_ = _3889_ & hart_id_i[16];
  assign _1329_ = _0051_ & _2950_;
  assign _1332_ = _2000_ & _2951_;
  assign _1335_ = _0473_ & _2952_;
  assign _1338_ = _0433_ & _2953_;
  assign _1341_ = _3743_ & _2954_;
  assign _1344_ = _3831_ & _2955_;
  assign _1347_ = _1994_ & _2956_;
  assign _1349_ = _0041_ & _0416_;
  assign _1352_ = _0029_ & _2957_;
  assign _1355_ = _0031_ & _2958_;
  assign _1358_ = _1996_ & _2959_;
  assign _1361_ = _0429_ & _2960_;
  assign _1364_ = _3893_ & _2961_;
  assign _1367_ = _0045_ & _2962_;
  assign _1370_ = _2004_ & _2963_;
  assign _1373_ = _0053_ & _2964_;
  assign _1375_ = _3889_ & hart_id_i[17];
  assign _1378_ = _0059_ & _2965_;
  assign _1381_ = _2006_ & _2966_;
  assign _1384_ = _0437_ & _2967_;
  assign _1387_ = _0439_ & _2968_;
  assign _1390_ = { _0021_, _0021_, _0021_ } & _2969_;
  assign _1393_ = { _3738_, _3738_, _3738_ } & _2970_;
  assign _1396_ = { _3741_, _3741_, _3741_ } & _2971_;
  assign _1399_ = { _2008_, _2008_, _2008_ } & _2972_;
  assign _1402_ = { _3831_, _3831_, _3831_ } & _2973_;
  assign _1405_ = { _0033_, _0033_, _0033_ } & _2974_;
  assign _1408_ = { _0041_, _0041_, _0041_ } & _2975_;
  assign _1411_ = { _2010_, _2010_, _2010_ } & _2976_;
  assign _1414_ = { _0475_, _0475_, _0475_ } & _2977_;
  assign _1417_ = { _0029_, _0029_, _0029_ } & _2978_;
  assign _1420_ = { _0039_, _0039_, _0039_ } & _2979_;
  assign _1423_ = { _0063_, _0063_, _0063_ } & _2980_;
  assign _1426_ = { _2012_, _2012_, _2012_ } & _2981_;
  assign _1429_ = { _3838_, _3838_, _3838_ } & _2982_;
  assign _1431_ = { _3889_, _3889_, _3889_ } & hart_id_i[2:0];
  assign _1433_ = { _3891_, _3891_, _3891_ } & _2983_;
  assign _1436_ = { _2000_, _2000_, _2000_ } & _2984_;
  assign _1439_ = { _0477_, _0477_, _0477_ } & _2985_;
  assign _1442_ = { _0479_, _0479_, _0479_ } & _2986_;
  assign _1444_ = _3743_ & _0417_;
  assign _1447_ = _3827_ & _2987_;
  assign _1450_ = _2024_ & _2988_;
  assign _1453_ = _3847_ & _2989_;
  assign _1456_ = _0033_ & _2990_;
  assign _1459_ = _2018_ & _2991_;
  assign _1462_ = _0481_ & _2992_;
  assign _1465_ = _0029_ & _2993_;
  assign _1468_ = _0063_ & _2994_;
  assign _1471_ = _2012_ & _2995_;
  assign _1474_ = _3838_ & _2996_;
  assign _1476_ = _3889_ & hart_id_i[12];
  assign _1479_ = _0059_ & _2997_;
  assign _1482_ = _2000_ & _2998_;
  assign _1485_ = _0469_ & _2999_;
  assign _1488_ = _0483_ & _3000_;
  assign _1490_ = _0159_ & debug_mode_i;
  assign _1492_ = _0157_ & _3001_;
  assign _1539_ = csr_restore_mret_i_t0 & _3003_;
  assign _1542_ = csr_restore_dret_i_t0 & _3004_;
  assign _1545_ = csr_save_cause_i_t0 & _3005_;
  assign _1547_ = nmi_mode_i_t0 & _0418_;
  assign _1550_ = { nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0 } & _3006_;
  assign _1552_ = nmi_mode_i_t0 & _0419_;
  assign _1555_ = { nmi_mode_i_t0, nmi_mode_i_t0 } & mstack_q[1:0];
  assign _1557_ = nmi_mode_i_t0 & _0420_;
  assign _1560_ = { csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0 } & _3007_;
  assign _1563_ = { csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0 } & _3008_;
  assign _1566_ = { csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0 } & _3009_;
  assign _1569_ = { nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0 } & _3010_;
  assign _1572_ = { debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0 } & _3011_;
  assign _1574_ = debug_mode_i_t0 & _0418_;
  assign _1577_ = { debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0 } & _3012_;
  assign _1579_ = debug_mode_i_t0 & _0419_;
  assign _1582_ = { debug_mode_i_t0, debug_mode_i_t0 } & _3013_;
  assign _1585_ = debug_mode_i_t0 & _3014_;
  assign _1587_ = debug_mode_i_t0 & _0421_;
  assign _1590_ = { debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0 } & _3015_;
  assign _1592_ = debug_mode_i_t0 & _0422_;
  assign _1594_ = debug_csr_save_i_t0 & _0423_;
  assign _1597_ = { debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0 } & _3012_;
  assign _1599_ = debug_csr_save_i_t0 & _0424_;
  assign _1602_ = { debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0 } & _3016_;
  assign _1605_ = { debug_csr_save_i_t0, debug_csr_save_i_t0 } & _3017_;
  assign _1607_ = debug_csr_save_i_t0 & _0072_;
  assign _1610_ = debug_csr_save_i_t0 & _3018_;
  assign _1613_ = { debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0 } & _3019_;
  assign _1616_ = debug_csr_save_i_t0 & _3020_;
  assign _1619_ = { debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0 } & _3021_;
  assign _1622_ = debug_csr_save_i_t0 & _3022_;
  assign _1625_ = { debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0 } & _3023_;
  assign _1628_ = debug_csr_save_i_t0 & _3024_;
  assign _1631_ = { debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0 } & _3025_;
  assign _1634_ = { csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0 } & _3026_;
  assign _1637_ = { csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0 } & _3027_;
  assign _1640_ = { csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0 } & _3028_;
  assign _1642_ = csr_save_cause_i_t0 & _0054_;
  assign _1645_ = csr_save_cause_i_t0 & _3029_;
  assign _1648_ = { csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0 } & _3030_;
  assign _1651_ = csr_save_cause_i_t0 & _3031_;
  assign _1654_ = { csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0 } & _3032_;
  assign _1657_ = { csr_save_cause_i_t0, csr_save_cause_i_t0 } & _3033_;
  assign _1660_ = csr_save_cause_i_t0 & _3034_;
  assign _1663_ = { csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0 } & _3035_;
  assign _1666_ = csr_restore_mret_i_t0 & _3036_;
  assign _1669_ = csr_restore_dret_i_t0 & _3037_;
  assign _1672_ = csr_save_cause_i_t0 & _3038_;
  assign _1675_ = { csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0 } & _3039_;
  assign _1678_ = { csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0 } & _3040_;
  assign _1681_ = { csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0 } & _3041_;
  assign _1684_ = csr_restore_mret_i_t0 & _3042_;
  assign _1687_ = csr_restore_dret_i_t0 & _3043_;
  assign _1690_ = csr_save_cause_i_t0 & _3044_;
  assign _1693_ = { csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0 } & _3045_;
  assign _1696_ = { csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0 } & _3046_;
  assign _1699_ = { csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0 } & _3047_;
  assign _1701_ = csr_restore_mret_i_t0 & _0421_;
  assign _1704_ = csr_restore_dret_i_t0 & _3048_;
  assign _1707_ = csr_save_cause_i_t0 & _3049_;
  assign _1709_ = debug_mode_i_t0 & _0010_[5];
  assign _1712_ = { csr_restore_mret_i_t0, csr_restore_mret_i_t0 } & _3050_;
  assign _1715_ = { csr_restore_dret_i_t0, csr_restore_dret_i_t0 } & _3051_;
  assign _1718_ = { csr_save_cause_i_t0, csr_save_cause_i_t0 } & _3052_;
  assign _1721_ = { _0025_, _0025_, _0025_, _0025_ } & _3053_;
  assign _1724_ = { _0059_, _0059_ } & _3054_;
  assign _1727_ = { _0059_, _0059_ } & _3055_;
  assign _1730_ = _0025_ & _3056_;
  assign _1732_ = _0025_ & dcsr_q[14];
  assign _1735_ = { _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_ } & dcsr_q[27:16];
  assign _1738_ = { _0059_, _0059_ } & _3057_;
  assign _1741_ = { _0025_, _0025_ } & _3058_;
  assign _1743_ = _0025_ & dcsr_q[5];
  assign _1745_ = _0025_ & dcsr_q[4];
  assign _1747_ = _0025_ & dcsr_q[3];
  assign _1750_ = _0025_ & _3059_;
  assign _1753_ = { _0025_, _0025_ } & _3060_;
  assign _1755_ = _0025_ & dcsr_q[11];
  assign _1758_ = { _3749_, _3749_ } & _3061_;
  assign _1760_ = _0025_ & dcsr_q[9];
  assign _1763_ = { _3747_, _3747_ } & _3062_;
  assign _1766_ = { _3827_, _3827_, _3827_, _3827_, _3827_, _3827_, _3827_, _3827_, _3827_, _3827_, _3827_, _3827_, _3827_, _3827_, _3827_, _3827_, _3827_, _3827_, _3827_, _3827_, _3827_, _3827_, _3827_, _3827_, _3827_, _3827_, _3827_, _3827_, _3827_, _3827_, _3827_, _3827_ } & _3063_;
  assign _1769_ = { _3831_, _3831_, _3831_, _3831_, _3831_, _3831_, _3831_, _3831_, _3831_, _3831_, _3831_, _3831_, _3831_, _3831_, _3831_, _3831_, _3831_, _3831_, _3831_, _3831_, _3831_, _3831_, _3831_, _3831_, _3831_, _3831_, _3831_, _3831_, _3831_, _3831_, _3831_, _3831_ } & _3063_;
  assign _1771_ = _0025_ & dcsr_q[10];
  assign _1773_ = _3838_ & _0425_;
  assign _1775_ = csr_we_int_t0 & _0020_;
  assign _1778_ = { csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0 } & _0048_;
  assign _1780_ = { csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0 } & _0046_;
  assign _1782_ = csr_we_int_t0 & _0040_;
  assign _1784_ = csr_we_int_t0 & _0032_;
  assign _1786_ = csr_we_int_t0 & _0030_;
  assign _1788_ = csr_we_int_t0 & _0028_;
  assign _1790_ = csr_we_int_t0 & _0024_;
  assign _1793_ = { csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0 } & _3064_;
  assign _1796_ = csr_we_int_t0 & _3065_;
  assign _1798_ = csr_we_int_t0 & _0062_;
  assign _1800_ = csr_we_int_t0 & _0038_;
  assign _1802_ = csr_we_int_t0 & _0044_;
  assign _1804_ = csr_we_int_t0 & _0052_;
  assign _1806_ = csr_we_int_t0 & _0050_;
  assign _1808_ = csr_we_int_t0 & _0058_;
  assign _1811_ = { csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0 } & _3066_;
  assign _1987_ = { csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0 } & _3067_;
  assign _1990_ = { mstatus_q_t0[1], mstatus_q_t0[1] } & _3050_;
  assign _1992_ = _3751_ & csr_wdata_int[0];
  assign _3242_ = _0727_ | _2071_;
  assign csr_wdata_int_t0 = _0730_ | _2074_;
  assign _3244_ = _0733_ | _2077_;
  assign _3246_ = _0736_ | _2080_;
  assign _3248_ = _0739_ | _2083_;
  assign _3250_ = _0741_ | _0740_;
  assign _3252_ = _0744_ | _2088_;
  assign _3254_ = _0747_ | _2091_;
  assign _3256_ = _0750_ | _2094_;
  assign _3258_ = _0753_ | _2097_;
  assign _3260_ = _0756_ | _2100_;
  assign _3262_ = _0759_ | _2103_;
  assign _3264_ = _0762_ | _2106_;
  assign _3266_ = _0764_ | _0763_;
  assign _3268_ = _0767_ | _2110_;
  assign _3270_ = _0770_ | _2113_;
  assign csr_rdata_o_t0[31] = _0773_ | _2116_;
  assign _3272_ = _0776_ | _2119_;
  assign _3274_ = _0779_ | _2122_;
  assign _3276_ = _0782_ | _2125_;
  assign _3278_ = _0785_ | _2128_;
  assign _3280_ = _0788_ | _2131_;
  assign _3282_ = _0791_ | _2134_;
  assign _3284_ = _0794_ | _2137_;
  assign _3286_ = _0797_ | _2140_;
  assign _3288_ = _0800_ | _2143_;
  assign _3290_ = _0803_ | _2146_;
  assign _3292_ = _0806_ | _2149_;
  assign _3294_ = _0809_ | _2152_;
  assign _3296_ = _0812_ | _2155_;
  assign _3298_ = _0815_ | _2158_;
  assign csr_rdata_o_t0[10:8] = _0818_ | _2161_;
  assign _3300_ = _0821_ | _2162_;
  assign _3302_ = _0824_ | _2163_;
  assign _3304_ = _0827_ | _2164_;
  assign _3306_ = _0830_ | _2165_;
  assign _3308_ = _0833_ | _2168_;
  assign _3310_ = _0836_ | _2169_;
  assign _3312_ = _0839_ | _2170_;
  assign _3314_ = _0842_ | _2171_;
  assign _3316_ = _0845_ | _2174_;
  assign _3318_ = _0848_ | _2177_;
  assign _3320_ = _0851_ | _2180_;
  assign _3322_ = _0854_ | _2183_;
  assign _3324_ = _0856_ | _0855_;
  assign _3326_ = _0859_ | _2186_;
  assign _3328_ = _0862_ | _2189_;
  assign _3330_ = _0865_ | _2192_;
  assign csr_rdata_o_t0[7] = _0868_ | _2195_;
  assign _3332_ = _0871_ | _2198_;
  assign _3334_ = _0874_ | _2201_;
  assign _3336_ = _0877_ | _2204_;
  assign _3338_ = _0880_ | _2205_;
  assign _3340_ = _0883_ | _2208_;
  assign _3342_ = _0886_ | _2209_;
  assign _3344_ = _0889_ | _2212_;
  assign _3346_ = _0892_ | _2215_;
  assign _3348_ = _0895_ | _2218_;
  assign _3350_ = _0898_ | _2221_;
  assign _3352_ = _0901_ | _2224_;
  assign _3354_ = _0904_ | _2225_;
  assign _3356_ = _0906_ | _2226_;
  assign _3358_ = _0909_ | _2227_;
  assign _3360_ = _0912_ | _2230_;
  assign _3362_ = _0915_ | _2233_;
  assign csr_rdata_o_t0[6:4] = _0918_ | _2236_;
  assign _3363_ = _0921_ | _2239_;
  assign _3365_ = _0924_ | _2242_;
  assign _3367_ = _0927_ | _2245_;
  assign _3369_ = _0930_ | _2248_;
  assign _3371_ = _0933_ | _2251_;
  assign _3373_ = _0936_ | _2254_;
  assign _3375_ = _0939_ | _2257_;
  assign _3377_ = _0942_ | _2260_;
  assign _3379_ = _0945_ | _2263_;
  assign _3381_ = _0948_ | _2266_;
  assign _3383_ = _0951_ | _2269_;
  assign _0019_ = _0954_ | _2272_;
  assign _3385_ = _0957_ | _2275_;
  assign _3387_ = _0960_ | _2278_;
  assign _3389_ = _0962_ | _0961_;
  assign _3391_ = _0965_ | _2282_;
  assign _3393_ = _0968_ | _2285_;
  assign _3395_ = _0971_ | _2286_;
  assign _3397_ = _0974_ | _2289_;
  assign _3399_ = _0977_ | _2292_;
  assign _3401_ = _0980_ | _2295_;
  assign _3403_ = _0983_ | _2296_;
  assign _3405_ = _0986_ | _2297_;
  assign _3407_ = _0989_ | _2300_;
  assign _3409_ = _0992_ | _2303_;
  assign _3411_ = _0995_ | _2304_;
  assign _3413_ = _0998_ | _2305_;
  assign _3415_ = _1000_ | _0999_;
  assign _3417_ = _1003_ | _2306_;
  assign _3419_ = _1006_ | _2309_;
  assign _3421_ = _1009_ | _2312_;
  assign csr_rdata_o_t0[3] = _1012_ | _2315_;
  assign _3423_ = _1015_ | _2316_;
  assign _3425_ = _1018_ | _2317_;
  assign _3427_ = _1021_ | _2318_;
  assign _3429_ = _1024_ | _2319_;
  assign _3431_ = _1027_ | _2320_;
  assign _3433_ = _1030_ | _2321_;
  assign _3435_ = _1033_ | _2322_;
  assign _3437_ = _1036_ | _2323_;
  assign _3439_ = _1039_ | _2324_;
  assign _3441_ = _1042_ | _2325_;
  assign _3443_ = _1045_ | _2326_;
  assign _3445_ = _1048_ | _2327_;
  assign _3447_ = _1050_ | _1049_;
  assign _3449_ = _1053_ | _2328_;
  assign _3451_ = _1056_ | _2329_;
  assign _3453_ = _1059_ | _2330_;
  assign csr_rdata_o_t0[11] = _1062_ | _2331_;
  assign _3455_ = _1065_ | _2332_;
  assign _3457_ = _1068_ | _2333_;
  assign _3459_ = _1071_ | _2334_;
  assign _3461_ = _1073_ | _1072_;
  assign _3463_ = _1076_ | _2335_;
  assign _3465_ = _1079_ | _2336_;
  assign _3467_ = _1082_ | _2337_;
  assign _3469_ = _1085_ | _2338_;
  assign _3471_ = _1088_ | _2339_;
  assign _3473_ = _1091_ | _2340_;
  assign _3475_ = _1094_ | _2341_;
  assign _3477_ = _1097_ | _2342_;
  assign _3479_ = _1099_ | _1098_;
  assign _3481_ = _1102_ | _2343_;
  assign _3483_ = _1105_ | _2344_;
  assign _3485_ = _1108_ | _2345_;
  assign csr_rdata_o_t0[21] = _1111_ | _2346_;
  assign _3486_ = _1114_ | _2349_;
  assign _3488_ = _1117_ | _2352_;
  assign _3490_ = _1120_ | _2355_;
  assign _3492_ = _1123_ | _2358_;
  assign _3494_ = _1126_ | _2361_;
  assign _3496_ = _1129_ | _2364_;
  assign _3498_ = _1132_ | _2367_;
  assign _3500_ = _1135_ | _2370_;
  assign _3502_ = _1138_ | _2373_;
  assign _3504_ = _1141_ | _2376_;
  assign _3506_ = _1144_ | _2379_;
  assign _0017_ = _1147_ | _2382_;
  assign _3508_ = _1150_ | _2385_;
  assign _3510_ = _1153_ | _2388_;
  assign _3512_ = _1156_ | _2391_;
  assign _3514_ = _1159_ | _2394_;
  assign _3516_ = _1162_ | _2397_;
  assign _3518_ = _1165_ | _2400_;
  assign _3520_ = _1168_ | _2403_;
  assign _3522_ = _1171_ | _2406_;
  assign _3524_ = _1174_ | _2409_;
  assign _3526_ = _1177_ | _2412_;
  assign _3528_ = _1180_ | _2415_;
  assign _3530_ = _1183_ | _2418_;
  assign _3532_ = _1186_ | _2421_;
  assign _3534_ = _1189_ | _2424_;
  assign _3536_ = _1192_ | _2427_;
  assign _3538_ = _1195_ | _2430_;
  assign _3540_ = _1198_ | _2433_;
  assign csr_rdata_o_t0[30:22] = _1201_ | _2436_;
  assign _3542_ = _1204_ | _2439_;
  assign _3544_ = _1207_ | _2440_;
  assign _3546_ = _1210_ | _2443_;
  assign _3548_ = _1213_ | _2444_;
  assign _3550_ = _1216_ | _2447_;
  assign _3552_ = _1219_ | _2450_;
  assign _3554_ = _1222_ | _2451_;
  assign _3556_ = _1225_ | _2452_;
  assign _3558_ = _1228_ | _2453_;
  assign _3560_ = _1231_ | _2456_;
  assign _3562_ = _1233_ | _2457_;
  assign _3564_ = _1236_ | _2460_;
  assign _3566_ = _1239_ | _2463_;
  assign csr_rdata_o_t0[15:13] = _1242_ | _2466_;
  assign _3568_ = _1245_ | _2467_;
  assign _3570_ = _1248_ | _2468_;
  assign _3572_ = _1251_ | _2469_;
  assign _3574_ = _1254_ | _2470_;
  assign _3576_ = _1257_ | _2471_;
  assign _3578_ = _1260_ | _2472_;
  assign _3580_ = _1263_ | _2473_;
  assign _3582_ = _1266_ | _2474_;
  assign _3584_ = _1269_ | _2477_;
  assign _3586_ = _1272_ | _2478_;
  assign _3588_ = _1275_ | _2481_;
  assign _3590_ = _1278_ | _2482_;
  assign _3592_ = _1280_ | _2483_;
  assign _3594_ = _1283_ | _2486_;
  assign _3596_ = _1286_ | _2489_;
  assign _3598_ = _1289_ | _2492_;
  assign csr_rdata_o_t0[20:18] = _1292_ | _2495_;
  assign _3600_ = _1295_ | _2496_;
  assign _3602_ = _1298_ | _2497_;
  assign _3604_ = _1301_ | _2498_;
  assign _3606_ = _1303_ | _1302_;
  assign _3608_ = _1306_ | _2499_;
  assign _3610_ = _1309_ | _2500_;
  assign _3612_ = _1312_ | _2501_;
  assign _3614_ = _1315_ | _2502_;
  assign _3616_ = _1318_ | _2503_;
  assign _3618_ = _1321_ | _2504_;
  assign _3620_ = _1324_ | _2505_;
  assign _3622_ = _1326_ | _1325_;
  assign _3624_ = _1329_ | _2508_;
  assign _3626_ = _1332_ | _2509_;
  assign _3628_ = _1335_ | _2512_;
  assign csr_rdata_o_t0[16] = _1338_ | _2513_;
  assign _3630_ = _1341_ | _2514_;
  assign _3632_ = _1344_ | _2515_;
  assign _3634_ = _1347_ | _2516_;
  assign _3636_ = _1349_ | _1348_;
  assign _3638_ = _1352_ | _2517_;
  assign _3640_ = _1355_ | _2518_;
  assign _3642_ = _1358_ | _2519_;
  assign _3644_ = _1361_ | _2520_;
  assign _3646_ = _1364_ | _2521_;
  assign _3648_ = _1367_ | _2522_;
  assign _3650_ = _1370_ | _2523_;
  assign _3652_ = _1373_ | _2524_;
  assign _3654_ = _1375_ | _1374_;
  assign _3656_ = _1378_ | _2525_;
  assign _3658_ = _1381_ | _2526_;
  assign _3660_ = _1384_ | _2527_;
  assign csr_rdata_o_t0[17] = _1387_ | _2528_;
  assign _3662_ = _1390_ | _2529_;
  assign _3664_ = _1393_ | _2532_;
  assign _3666_ = _1396_ | _2533_;
  assign _3668_ = _1399_ | _2534_;
  assign _3670_ = _1402_ | _2535_;
  assign _3672_ = _1405_ | _2536_;
  assign _3674_ = _1408_ | _2537_;
  assign _3676_ = _1411_ | _2538_;
  assign _3678_ = _1414_ | _2541_;
  assign _3680_ = _1417_ | _2542_;
  assign _3682_ = _1420_ | _2545_;
  assign _3684_ = _1423_ | _2546_;
  assign _3686_ = _1426_ | _2547_;
  assign _3688_ = _1429_ | _2548_;
  assign _3690_ = _1431_ | _2549_;
  assign _3692_ = _1433_ | _2550_;
  assign _3694_ = _1436_ | _2551_;
  assign _3696_ = _1439_ | _2554_;
  assign csr_rdata_o_t0[2:0] = _1442_ | _2557_;
  assign _3698_ = _1444_ | _1443_;
  assign _3700_ = _1447_ | _2558_;
  assign _3702_ = _1450_ | _2561_;
  assign _3704_ = _1453_ | _2562_;
  assign _3706_ = _1456_ | _2563_;
  assign _3708_ = _1459_ | _2564_;
  assign _3710_ = _1462_ | _2567_;
  assign _3712_ = _1465_ | _2568_;
  assign _3714_ = _1468_ | _2569_;
  assign _3716_ = _1471_ | _2572_;
  assign _3718_ = _1474_ | _2573_;
  assign _3720_ = _1476_ | _1475_;
  assign _3722_ = _1479_ | _2574_;
  assign _3724_ = _1482_ | _2575_;
  assign _3726_ = _1485_ | _2578_;
  assign csr_rdata_o_t0[12] = _1488_ | _2581_;
  assign _3727_ = _1490_ | _1489_;
  assign illegal_csr_t0 = _1492_ | _1491_;
  assign _3787_ = _1539_ | _2603_;
  assign _3789_ = _1542_ | _2606_;
  assign mstatus_d_t0[5] = _1545_ | _2609_;
  assign _0106_ = _1547_ | _1546_;
  assign _0086_ = _1550_ | _2614_;
  assign _0108_ = _1552_ | _1551_;
  assign _0114_[1:0] = _1555_ | _2617_;
  assign _0114_[2] = _1557_ | _1556_;
  assign _3791_ = _1560_ | _2620_;
  assign _3793_ = _1563_ | _2623_;
  assign mstatus_d_t0[4:2] = _1566_ | _2626_;
  assign _0082_ = _1569_ | _2629_;
  assign _0069_ = _1572_ | _2632_;
  assign _0094_ = _1574_ | _1573_;
  assign _0071_ = _1577_ | _2637_;
  assign _0096_ = _1579_ | _1578_;
  assign _0110_[1:0] = _1582_ | _2640_;
  assign _0110_[2] = _1585_ | _2641_;
  assign _0100_ = _1587_ | _1586_;
  assign _0076_ = _1590_ | _2642_;
  assign _0102_ = _1592_ | _1591_;
  assign _0080_ = _1594_ | _1593_;
  assign _0027_ = _1597_ | _2647_;
  assign _0078_ = _1599_ | _1598_;
  assign _0112_ = _1602_ | _2650_;
  assign _0104_ = _1605_ | _2653_;
  assign _0055_ = _1607_ | _1606_;
  assign _0092_ = _1610_ | _2654_;
  assign _0061_ = _1613_ | _2655_;
  assign _0084_ = _1616_ | _2656_;
  assign _0037_ = _1619_ | _2659_;
  assign _0088_ = _1622_ | _2660_;
  assign _0043_ = _1625_ | _2661_;
  assign _0090_ = _1628_ | _2662_;
  assign _0098_ = _1631_ | _2665_;
  assign _3795_ = _1634_ | _2668_;
  assign _3797_ = _1637_ | _2671_;
  assign _0035_ = _1640_ | _2674_;
  assign mstack_en_t0 = _1642_ | _1641_;
  assign depc_en_t0 = _1645_ | _2675_;
  assign depc_d_t0 = _1648_ | _2678_;
  assign dcsr_en_t0 = _1651_ | _2679_;
  assign dcsr_d_t0[8:6] = _1654_ | _2680_;
  assign dcsr_d_t0[1:0] = _1657_ | _2683_;
  assign mtval_en_t0 = _1660_ | _2684_;
  assign mtval_d_t0 = _1663_ | _2685_;
  assign _3799_ = _1666_ | _2686_;
  assign _3801_ = _1669_ | _2687_;
  assign mcause_en_t0 = _1672_ | _2688_;
  assign _3803_ = _1675_ | _2691_;
  assign _3805_ = _1678_ | _2694_;
  assign mcause_d_t0 = _1681_ | _2697_;
  assign _3807_ = _1684_ | _2698_;
  assign _3809_ = _1687_ | _2699_;
  assign mepc_en_t0 = _1690_ | _2700_;
  assign _3811_ = _1693_ | _2703_;
  assign _3813_ = _1696_ | _2706_;
  assign mepc_d_t0 = _1699_ | _2707_;
  assign _3815_ = _1701_ | _1700_;
  assign _3817_ = _1704_ | _2708_;
  assign mstatus_en_t0 = _1707_ | _2709_;
  assign _0110_[3] = _1709_ | _1708_;
  assign _3819_ = _1712_ | _2712_;
  assign _3821_ = _1715_ | _2715_;
  assign priv_mode_if_o_t0 = _1718_ | _2716_;
  assign _0023_[31:28] = _1721_ | _2719_;
  assign _0057_[5:4] = _1724_ | _2722_;
  assign _0057_[3:2] = _1727_ | _2723_;
  assign _0023_[15] = _1730_ | _2724_;
  assign _0023_[14] = _1732_ | _1731_;
  assign _0023_[27:16] = _1735_ | _2727_;
  assign _0057_[1:0] = _1738_ | _2728_;
  assign _0023_[1:0] = _1741_ | _2731_;
  assign _0023_[5] = _1743_ | _1742_;
  assign _0023_[4] = _1745_ | _1744_;
  assign _0023_[3] = _1747_ | _1746_;
  assign _0023_[2] = _1750_ | _2732_;
  assign _0023_[13:12] = _1753_ | _2733_;
  assign _0023_[11] = _1755_ | _1754_;
  assign _0067_ = _1758_ | _2736_;
  assign _0023_[9] = _1760_ | _1759_;
  assign _0074_ = _1763_ | _2739_;
  assign _0049_ = _1766_ | _2742_;
  assign _0047_ = _1769_ | _2745_;
  assign _0023_[10] = _1771_ | _1770_;
  assign _0065_ = _1773_ | _1772_;
  assign cpuctrl_we_t0 = _1775_ | _1774_;
  assign mhpmcounterh_we_t0 = _1778_ | _2750_;
  assign mhpmcounter_we_t0 = _1780_ | _2751_;
  assign mcountinhibit_we_t0 = _1782_ | _1781_;
  assign dscratch1_en_t0 = _1784_ | _1783_;
  assign dscratch0_en_t0 = _1786_ | _1785_;
  assign _0005_ = _1788_ | _1787_;
  assign _0003_ = _1790_ | _1789_;
  assign { dcsr_d_t0[31:9], _0001_[8:6], dcsr_d_t0[5:2], _0001_[1:0] } = _1793_ | _2752_;
  assign mtvec_en_t0 = _1796_ | _2753_;
  assign _0015_ = _1798_ | _1797_;
  assign _0007_ = _1800_ | _1799_;
  assign _0009_ = _1802_ | _1801_;
  assign mscratch_en_t0 = _1804_ | _1803_;
  assign mie_en_t0 = _1806_ | _1805_;
  assign _0013_ = _1808_ | _1807_;
  assign { _0011_[5:2], mstatus_d_t0[1:0] } = _1811_ | _2756_;
  assign mtvec_d_t0 = _1987_ | _2759_;
  assign priv_mode_lsu_o_t0 = _1990_ | _2762_;
  assign \gen_trigger_regs.tselect_d_t0  = _1992_ | _1991_;
  assign _0346_ = ~ { 27'h0000000, csr_addr_i_t0[4:0] };
  assign _1516_ = { 27'h0000000, csr_addr_i[4:0] } & _0346_;
  assign _2594_ = { 27'h0000000, csr_addr_i[4:0] } | { 27'h0000000, csr_addr_i_t0[4:0] };
  assign _0426_ = - _1516_;
  assign _0427_ = - _2594_;
  assign _3002_ = _0426_ ^ _0427_;
  assign _3761_ = _3002_ | { 27'h0000000, csr_addr_i_t0[4:0] };
  assign _0412_ = ~ dscratch1_q[31];
  assign _0413_ = ~ _3386_;
  assign _0414_ = ~ dscratch1_q[21];
  assign _0415_ = ~ dscratch1_q[16];
  assign _0416_ = ~ dscratch1_q[17];
  assign _0417_ = ~ \gen_trigger_regs.selected_tmatch_value [12];
  assign _0420_ = ~ mstack_q[2];
  assign _0418_ = ~ _0006_;
  assign _0419_ = ~ _0008_;
  assign _0422_ = ~ _0014_;
  assign _0423_ = ~ _0004_;
  assign _0424_ = ~ _0002_;
  assign _0421_ = ~ _0012_;
  assign _0425_ = ~ csr_mtvec_init_i;
  assign _0156_ = | { _3964_, _3962_, _3960_, _3958_, _3956_, _3892_, _3890_, _3888_, _3886_, _3884_, _3882_, _3880_, _3878_, _3876_, _3874_, _3872_, _3870_, _3868_, _3866_, _3864_, _3862_, _3860_, _3858_, _3856_, _3854_, _3852_, _3850_, _3848_, _3844_, _3843_, _3842_, _3841_, _3840_, _3839_, _3837_, _3833_, _3832_, _3828_, _3824_, _3823_, _3742_, _3740_, _3737_ };
  assign _0158_ = | { _3836_, _3835_, _3834_, _3822_ };
  assign _0154_ = | { _3954_, _3930_, _3928_, _3926_, _3924_, _3922_, _3920_, _3918_, _3916_, _3914_, _3912_, _3910_, _3908_, _3906_, _3904_, _3902_, _3900_, _3898_, _3896_, _3894_ };
  assign _0160_ = | { _3735_, _3784_ };
  assign _0162_ = | { _3890_, _3740_ };
  assign _0172_ = ~ _3890_;
  assign _0176_ = ~ _3950_;
  assign _0188_ = ~ _0162_;
  assign _0347_ = ~ _0115_;
  assign _0349_ = ~ illegal_csr;
  assign _0351_ = ~ _3776_;
  assign _0353_ = ~ csr_wdata_i;
  assign _0355_ = ~ mstatus_err;
  assign _0357_ = ~ _3782_;
  assign _0177_ = ~ _3948_;
  assign _0348_ = ~ _3966_;
  assign _0350_ = ~ illegal_csr_write;
  assign _0352_ = ~ illegal_csr_priv;
  assign _0354_ = ~ csr_rdata_o;
  assign _0356_ = ~ mtvec_err;
  assign _0358_ = ~ cpuctrl_err;
  assign _0649_ = _0063_ & _0171_;
  assign _0652_ = _3891_ & _0173_;
  assign _0655_ = _3838_ & _0175_;
  assign _0658_ = _3951_ & _0177_;
  assign _0661_ = _3741_ & _0179_;
  assign _0664_ = _3893_ & _0171_;
  assign _0667_ = _3827_ & _0179_;
  assign _0670_ = _0033_ & _0183_;
  assign _0673_ = _0063_ & _0180_;
  assign _0676_ = _0051_ & _0173_;
  assign _0679_ = _3743_ & _0185_;
  assign _0682_ = _3847_ & _0187_;
  assign _0685_ = _0163_ & _0179_;
  assign _0688_ = _0041_ & _0186_;
  assign _0691_ = _0025_ & _0189_;
  assign _0694_ = _0053_ & _0174_;
  assign _1517_ = _0116_ & _0348_;
  assign _1520_ = illegal_csr_t0 & _0350_;
  assign _1523_ = _3777_ & _0352_;
  assign _1526_ = csr_wdata_i_t0 & _0354_;
  assign _1527_ = mstatus_err_t0 & _0356_;
  assign _1530_ = _3783_ & _0358_;
  assign _0650_ = _0025_ & _0170_;
  assign _0653_ = _0053_ & _0172_;
  assign _0656_ = _0045_ & _0174_;
  assign _0659_ = _3949_ & _0176_;
  assign _0662_ = _3743_ & _0178_;
  assign _0665_ = _0025_ & _0180_;
  assign _0668_ = _3743_ & _0181_;
  assign _0671_ = _0041_ & _0182_;
  assign _0674_ = _3893_ & _0170_;
  assign _0677_ = _0053_ & _0184_;
  assign _0680_ = _0021_ & _0179_;
  assign _0683_ = _3831_ & _0186_;
  assign _0686_ = _3743_ & _0188_;
  assign _0689_ = _3847_ & _0183_;
  assign _0692_ = _0029_ & _0171_;
  assign _0695_ = _3838_ & _0173_;
  assign _1518_ = _3762_ & _0347_;
  assign _1521_ = illegal_csr_write_t0 & _0349_;
  assign _1524_ = illegal_csr_priv_t0 & _0351_;
  assign _0576_ = csr_rdata_o_t0 & _0353_;
  assign _1528_ = mtvec_err_t0 & _0355_;
  assign _1531_ = cpuctrl_err_t0 & _0357_;
  assign _0651_ = _0063_ & _0025_;
  assign _0654_ = _3891_ & _0053_;
  assign _0657_ = _3838_ & _0045_;
  assign _0660_ = _3951_ & _3949_;
  assign _0663_ = _3741_ & _3743_;
  assign _0666_ = _3893_ & _0025_;
  assign _0669_ = _3827_ & _3743_;
  assign _0672_ = _0033_ & _0041_;
  assign _0675_ = _0063_ & _3893_;
  assign _0678_ = _0051_ & _0053_;
  assign _0681_ = _3743_ & _0021_;
  assign _0684_ = _3847_ & _3831_;
  assign _0687_ = _0163_ & _3743_;
  assign _0690_ = _0041_ & _3847_;
  assign _0693_ = _0025_ & _0029_;
  assign _0696_ = _0053_ & _3838_;
  assign _1519_ = _0116_ & _3762_;
  assign _1522_ = illegal_csr_t0 & illegal_csr_write_t0;
  assign _1525_ = _3777_ & illegal_csr_priv_t0;
  assign _0577_ = csr_wdata_i_t0 & csr_rdata_o_t0;
  assign _1529_ = mstatus_err_t0 & mtvec_err_t0;
  assign _1532_ = _3783_ & cpuctrl_err_t0;
  assign _2053_ = _0649_ | _0650_;
  assign _2054_ = _0652_ | _0653_;
  assign _2055_ = _0655_ | _0656_;
  assign _2056_ = _0658_ | _0659_;
  assign _2057_ = _0661_ | _0662_;
  assign _2058_ = _0664_ | _0665_;
  assign _2059_ = _0667_ | _0668_;
  assign _2060_ = _0670_ | _0671_;
  assign _2061_ = _0673_ | _0674_;
  assign _2062_ = _0676_ | _0677_;
  assign _2063_ = _0679_ | _0680_;
  assign _2064_ = _0682_ | _0683_;
  assign _2065_ = _0685_ | _0686_;
  assign _2066_ = _0688_ | _0689_;
  assign _2067_ = _0691_ | _0692_;
  assign _2068_ = _0694_ | _0695_;
  assign _2595_ = _1517_ | _1518_;
  assign _2596_ = _1520_ | _1521_;
  assign _2597_ = _1523_ | _1524_;
  assign _2598_ = _1526_ | _0576_;
  assign _2599_ = _1527_ | _1528_;
  assign _2600_ = _1530_ | _1531_;
  assign _1998_ = _2053_ | _0651_;
  assign _2002_ = _2054_ | _0654_;
  assign _2014_ = _2055_ | _0657_;
  assign _2016_ = _2056_ | _0660_;
  assign _2022_ = _2057_ | _0663_;
  assign _2020_ = _2058_ | _0666_;
  assign _1994_ = _2059_ | _0669_;
  assign _1996_ = _2060_ | _0672_;
  assign _2004_ = _2061_ | _0675_;
  assign _2006_ = _2062_ | _0678_;
  assign _2008_ = _2063_ | _0681_;
  assign _2010_ = _2064_ | _0684_;
  assign _2024_ = _2065_ | _0687_;
  assign _2018_ = _2066_ | _0690_;
  assign _2012_ = _2067_ | _0693_;
  assign _2000_ = _2068_ | _0696_;
  assign _3775_ = _2595_ | _1519_;
  assign _3777_ = _2596_ | _1522_;
  assign _3779_ = _2597_ | _1525_;
  assign _3781_ = _2598_ | _0577_;
  assign _3783_ = _2599_ | _1529_;
  assign csr_shadow_err_o_t0 = _2600_ | _1532_;
  assign _1997_ = _3839_ | _3822_;
  assign _2001_ = _3890_ | _3842_;
  assign _2013_ = _3837_ | _3841_;
  assign _2015_ = _3950_ | _3948_;
  assign _2021_ = _3740_ | _3742_;
  assign _2019_ = _3892_ | _3822_;
  assign _1993_ = _3826_ | _3742_;
  assign _1995_ = _3834_ | _3833_;
  assign _2003_ = _3839_ | _3892_;
  assign _2005_ = _3843_ | _3842_;
  assign _2007_ = _3742_ | _3832_;
  assign _2009_ = _3846_ | _3830_;
  assign _2023_ = _0162_ | _3742_;
  assign _2017_ = _3833_ | _3846_;
  assign _2011_ = _3822_ | _3836_;
  assign _1999_ = _3842_ | _3837_;
  assign _0430_ = | { _1997_, _3841_, _3840_ };
  assign _0434_ = | { _1997_, _3841_, _3837_ };
  assign _0440_ = | { _3824_, _2007_, _3740_ };
  assign _0442_ = | { _3840_, _3839_, _2011_ };
  assign _0444_ = | { _3835_, _3834_, _3833_, _3824_, _2007_, _2009_, _3740_ };
  assign _0452_ = | { _3828_, _3824_, _2007_, _3740_ };
  assign _0454_ = | { _3843_, _3842_, _3837_ };
  assign _0456_ = | { _3841_, _3840_, _3839_, _2019_ };
  assign _0458_ = | { _3836_, _3835_, _3834_, _3828_, _3824_, _2007_, _3740_, _2017_ };
  assign _0446_ = | { _3954_, _3934_, _3932_, _3930_, _3928_, _3926_, _3924_, _3922_, _3920_, _3918_, _3916_, _3914_, _3912_, _3910_, _3908_, _3906_, _3904_, _3902_, _3900_, _3898_, _3896_, _3894_ };
  assign _0448_ = | { _3946_, _3944_, _3942_ };
  assign _0450_ = | { _3954_, _3940_, _3938_, _3936_, _3934_, _3932_, _3930_, _3928_, _3926_, _3924_, _3922_, _3920_, _3918_, _3916_, _3914_, _3912_, _3910_, _3908_, _3906_, _3904_, _3902_, _3900_, _3898_, _3896_, _3894_ };
  assign _0460_ = | { _2021_, _3828_, _3824_ };
  assign _0462_ = | { _3841_, _3839_, _3837_, _2019_ };
  assign _0464_ = | { _2021_, _3836_, _3835_, _3834_, _3828_, _3824_, _2017_ };
  assign _0466_ = | { _3828_, _3824_, _3742_ };
  assign _0470_ = | { _3835_, _3834_, _3828_, _3824_, _3742_, _2017_ };
  assign _0438_ = | { _1995_, _1993_, _3844_, _3836_, _3835_, _3828_, _3822_ };
  assign _0472_ = | { _3841_, _3839_, _2019_ };
  assign _0432_ = | { _1995_, _1993_, _3844_, _3836_, _3835_, _3828_ };
  assign _0428_ = | { _1993_, _3844_, _3828_ };
  assign _0436_ = | { _2003_, _3841_, _3837_ };
  assign _0474_ = | { _3824_, _2007_, _3740_, _3737_ };
  assign _0476_ = | { _3841_, _3840_, _3839_, _2011_ };
  assign _0478_ = | { _3835_, _3834_, _3833_, _3824_, _2007_, _2009_, _3740_, _3737_ };
  assign _0480_ = | { _3828_, _3824_, _2023_ };
  assign _0468_ = | { _3841_, _3839_, _2011_ };
  assign _0482_ = | { _3835_, _3834_, _3828_, _3824_, _2017_, _2023_ };
  assign _3241_ = _3731_ ? _0117_ : _3780_;
  assign csr_wdata_int = _0160_ ? csr_wdata_i : _3241_;
  assign _3243_ = _3742_ ? \gen_trigger_regs.selected_tmatch_value [31] : _0016_[63];
  assign _3245_ = _3830_ ? _0016_[31] : _0018_[31];
  assign _3247_ = _1993_ ? _3243_ : _3245_;
  assign _3249_ = _3833_ ? 1'h1 : dscratch1_q[31];
  assign _3251_ = _3835_ ? dscratch0_q[31] : csr_depc_o[31];
  assign _3253_ = _1995_ ? _3249_ : _3251_;
  assign _3255_ = _0428_ ? _3247_ : _3253_;
  assign _3257_ = _3822_ ? dcsr_q[31] : mtval_q[31];
  assign _3259_ = _3840_ ? mcause_q[5] : csr_mepc_o[31];
  assign _3261_ = _1997_ ? _3257_ : _3259_;
  assign _3263_ = _3837_ ? csr_mtvec_o[31] : mscratch_q[31];
  assign _3265_ = _3888_ ? hart_id_i[31] : 1'h0;
  assign _3267_ = _1999_ ? _3263_ : _3265_;
  assign _3269_ = _0430_ ? _3261_ : _3267_;
  assign csr_rdata_o[31] = _0432_ ? _3255_ : _3269_;
  assign _3271_ = _3742_ ? \gen_trigger_regs.selected_tmatch_value [10:8] : _0016_[42:40];
  assign _3273_ = _3830_ ? _0016_[10:8] : _0018_[10:8];
  assign _3275_ = _1993_ ? _3271_ : _3273_;
  assign _3277_ = _3833_ ? mcountinhibit[10:8] : dscratch1_q[10:8];
  assign _3279_ = _3835_ ? dscratch0_q[10:8] : csr_depc_o[10:8];
  assign _3281_ = _1995_ ? _3277_ : _3279_;
  assign _3283_ = _0428_ ? _3275_ : _3281_;
  assign _3285_ = _3822_ ? dcsr_q[10:8] : mtval_q[10:8];
  assign _3287_ = _3841_ ? csr_mepc_o[10:8] : csr_mtvec_o[10:8];
  assign _3289_ = _1997_ ? _3285_ : _3287_;
  assign _3291_ = _3842_ ? mscratch_q[10:8] : 3'h1;
  assign _3293_ = _3888_ ? hart_id_i[10:8] : 3'h0;
  assign _3295_ = _2001_ ? _3291_ : _3293_;
  assign _3297_ = _0434_ ? _3289_ : _3295_;
  assign csr_rdata_o[10:8] = _0432_ ? _3283_ : _3297_;
  assign _3299_ = _3742_ ? \gen_trigger_regs.selected_tmatch_value [7] : _0016_[39];
  assign _3301_ = _3830_ ? _0016_[7] : _0018_[7];
  assign _3303_ = _1993_ ? _3299_ : _3301_;
  assign _3305_ = _3833_ ? mcountinhibit[7] : dscratch1_q[7];
  assign _3307_ = _3836_ ? csr_depc_o[7] : dcsr_q[7];
  assign _3309_ = _3835_ ? dscratch0_q[7] : _3307_;
  assign _3311_ = _1995_ ? _3305_ : _3309_;
  assign _3313_ = _0428_ ? _3303_ : _3311_;
  assign _3315_ = _3892_ ? irq_timer_i : mtval_q[7];
  assign _3317_ = _3841_ ? csr_mepc_o[7] : csr_mtvec_o[7];
  assign _3319_ = _2003_ ? _3315_ : _3317_;
  assign _3321_ = _3842_ ? mscratch_q[7] : mie_q[16];
  assign _3323_ = _3888_ ? hart_id_i[7] : 1'h0;
  assign _3325_ = _3823_ ? mstatus_q[4] : _3323_;
  assign _3327_ = _2005_ ? _3321_ : _3325_;
  assign _3329_ = _0436_ ? _3319_ : _3327_;
  assign csr_rdata_o[7] = _0438_ ? _3313_ : _3329_;
  assign _3331_ = _3832_ ? { 1'h0, cpuctrl_q[5:4] } : \gen_trigger_regs.selected_tmatch_value [6:4];
  assign _3333_ = _3740_ ? 3'h4 : _0016_[38:36];
  assign _3335_ = _2007_ ? _3331_ : _3333_;
  assign _3337_ = _3830_ ? _0016_[6:4] : _0018_[6:4];
  assign _3339_ = _3834_ ? dscratch1_q[6:4] : dscratch0_q[6:4];
  assign _3341_ = _3833_ ? mcountinhibit[6:4] : _3339_;
  assign _3343_ = _2009_ ? _3337_ : _3341_;
  assign _3345_ = _0440_ ? _3335_ : _3343_;
  assign _3347_ = _3836_ ? csr_depc_o[6:4] : dcsr_q[6:4];
  assign _3349_ = _3839_ ? mtval_q[6:4] : { 2'h0, mcause_q[4] };
  assign _3351_ = _2011_ ? _3347_ : _3349_;
  assign _3353_ = _3841_ ? csr_mepc_o[6:4] : csr_mtvec_o[6:4];
  assign _3355_ = _3888_ ? hart_id_i[6:4] : 3'h0;
  assign _3357_ = _3842_ ? mscratch_q[6:4] : _3355_;
  assign _3359_ = _2013_ ? _3353_ : _3357_;
  assign _3361_ = _0442_ ? _3351_ : _3359_;
  assign csr_rdata_o[6:4] = _0444_ ? _3345_ : _3361_;
  assign _2826_ = _3932_ ? 32'd4096 : 32'd2048;
  assign _3364_ = _0154_ ? 32'd0 : _2826_;
  assign _3366_ = _3938_ ? 32'd512 : 32'd256;
  assign _3368_ = _3936_ ? 32'd1024 : _3366_;
  assign _3370_ = _0446_ ? _3364_ : _3368_;
  assign _3372_ = _3944_ ? 32'd64 : 32'd32;
  assign _3374_ = _3942_ ? 32'd128 : _3372_;
  assign _3376_ = _3948_ ? 32'd16 : 32'd8;
  assign _3378_ = _3952_ ? 32'd4 : 32'd1;
  assign _3380_ = _2015_ ? _3376_ : _3378_;
  assign _3382_ = _0448_ ? _3374_ : _3380_;
  assign _0018_ = _0450_ ? _3370_ : _3382_;
  assign _3384_ = _3832_ ? cpuctrl_q[3] : \gen_trigger_regs.selected_tmatch_value [3];
  assign _3386_ = _3826_ ? _0016_[35] : _0016_[3];
  assign _3388_ = _3740_ ? 1'h1 : _3386_;
  assign _3390_ = _2007_ ? _3384_ : _3388_;
  assign _3392_ = _3846_ ? _0018_[3] : mcountinhibit[3];
  assign _3394_ = _3835_ ? dscratch0_q[3] : csr_depc_o[3];
  assign _3396_ = _3834_ ? dscratch1_q[3] : _3394_;
  assign _3398_ = _2017_ ? _3392_ : _3396_;
  assign _3400_ = _0452_ ? _3390_ : _3398_;
  assign _3402_ = _3822_ ? dcsr_q[3] : irq_software_i;
  assign _3404_ = _3840_ ? mcause_q[3] : csr_mepc_o[3];
  assign _3406_ = _3839_ ? mtval_q[3] : _3404_;
  assign _3408_ = _2019_ ? _3402_ : _3406_;
  assign _3410_ = _3842_ ? mscratch_q[3] : mie_q[17];
  assign _3412_ = _3837_ ? csr_mtvec_o[3] : _3410_;
  assign _3414_ = _3888_ ? hart_id_i[3] : 1'h0;
  assign _3416_ = _3823_ ? mstatus_q[5] : _3414_;
  assign _3418_ = _0454_ ? _3412_ : _3416_;
  assign _3420_ = _0456_ ? _3408_ : _3418_;
  assign csr_rdata_o[3] = _0458_ ? _3400_ : _3420_;
  assign _3422_ = _3742_ ? \gen_trigger_regs.selected_tmatch_value [11] : _0016_[43];
  assign _3424_ = _3830_ ? _0016_[11] : _0018_[11];
  assign _3426_ = _1993_ ? _3422_ : _3424_;
  assign _3428_ = _3833_ ? mcountinhibit[11] : dscratch1_q[11];
  assign _3430_ = _3836_ ? csr_depc_o[11] : dcsr_q[11];
  assign _3432_ = _3835_ ? dscratch0_q[11] : _3430_;
  assign _3434_ = _1995_ ? _3428_ : _3432_;
  assign _3436_ = _0428_ ? _3426_ : _3434_;
  assign _3438_ = _3892_ ? irq_external_i : mtval_q[11];
  assign _3440_ = _3841_ ? csr_mepc_o[11] : csr_mtvec_o[11];
  assign _3442_ = _2003_ ? _3438_ : _3440_;
  assign _3444_ = _3842_ ? mscratch_q[11] : mie_q[15];
  assign _3446_ = _3888_ ? hart_id_i[11] : 1'h0;
  assign _3448_ = _3823_ ? mstatus_q[2] : _3446_;
  assign _3450_ = _2005_ ? _3444_ : _3448_;
  assign _3452_ = _0436_ ? _3442_ : _3450_;
  assign csr_rdata_o[11] = _0438_ ? _3436_ : _3452_;
  assign _3454_ = _3742_ ? \gen_trigger_regs.selected_tmatch_value [21] : _0016_[53];
  assign _3456_ = _3830_ ? _0016_[21] : _0018_[21];
  assign _3458_ = _1993_ ? _3454_ : _3456_;
  assign _3460_ = _3833_ ? 1'h1 : dscratch1_q[21];
  assign _3462_ = _3836_ ? csr_depc_o[21] : dcsr_q[21];
  assign _3464_ = _3835_ ? dscratch0_q[21] : _3462_;
  assign _3466_ = _1995_ ? _3460_ : _3464_;
  assign _3468_ = _0428_ ? _3458_ : _3466_;
  assign _3470_ = _3892_ ? irq_fast_i[5] : mtval_q[21];
  assign _3472_ = _3841_ ? csr_mepc_o[21] : csr_mtvec_o[21];
  assign _3474_ = _2003_ ? _3470_ : _3472_;
  assign _3476_ = _3842_ ? mscratch_q[21] : mie_q[5];
  assign _3478_ = _3888_ ? hart_id_i[21] : 1'h0;
  assign _3480_ = _3823_ ? mstatus_q[0] : _3478_;
  assign _3482_ = _2005_ ? _3476_ : _3480_;
  assign _3484_ = _0436_ ? _3474_ : _3482_;
  assign csr_rdata_o[21] = _0438_ ? _3468_ : _3484_;
  assign _2883_ = _3932_ ? \mhpmcounter[12]  : \mhpmcounter[11] ;
  assign _3487_ = _0154_ ? 64'h0000000000000000 : _2883_;
  assign _3489_ = _3938_ ? \mhpmcounter[9]  : \mhpmcounter[8] ;
  assign _3491_ = _3936_ ? \mhpmcounter[10]  : _3489_;
  assign _3493_ = _0446_ ? _3487_ : _3491_;
  assign _3495_ = _3944_ ? \mhpmcounter[6]  : \mhpmcounter[5] ;
  assign _3497_ = _3942_ ? \mhpmcounter[7]  : _3495_;
  assign _3499_ = _3948_ ? \mhpmcounter[4]  : \mhpmcounter[3] ;
  assign _3501_ = _3952_ ? \mhpmcounter[2]  : \mhpmcounter[0] ;
  assign _3503_ = _2015_ ? _3499_ : _3501_;
  assign _3505_ = _0448_ ? _3497_ : _3503_;
  assign _0016_ = _0450_ ? _3493_ : _3505_;
  assign _3507_ = _3742_ ? \gen_trigger_regs.selected_tmatch_value [30:22] : 9'h0a0;
  assign _3509_ = _3826_ ? _0016_[62:54] : _0016_[30:22];
  assign _3511_ = _2021_ ? _3507_ : _3509_;
  assign _3513_ = _3846_ ? _0018_[30:22] : 9'h1ff;
  assign _3515_ = _3835_ ? dscratch0_q[30:22] : csr_depc_o[30:22];
  assign _3517_ = _3834_ ? dscratch1_q[30:22] : _3515_;
  assign _3519_ = _2017_ ? _3513_ : _3517_;
  assign _3521_ = _0460_ ? _3511_ : _3519_;
  assign _3523_ = _3822_ ? dcsr_q[30:22] : irq_fast_i[14:6];
  assign _3525_ = _3841_ ? csr_mepc_o[30:22] : csr_mtvec_o[30:22];
  assign _3527_ = _3839_ ? mtval_q[30:22] : _3525_;
  assign _3529_ = _2019_ ? _3523_ : _3527_;
  assign _3531_ = _3842_ ? mscratch_q[30:22] : mie_q[14:6];
  assign _3533_ = _3888_ ? hart_id_i[30:22] : 9'h000;
  assign _3535_ = _3890_ ? 9'h100 : _3533_;
  assign _3537_ = _2005_ ? _3531_ : _3535_;
  assign _3539_ = _0462_ ? _3529_ : _3537_;
  assign csr_rdata_o[30:22] = _0464_ ? _3521_ : _3539_;
  assign _3541_ = _3826_ ? _0016_[47:45] : _0016_[15:13];
  assign _3543_ = _3742_ ? \gen_trigger_regs.selected_tmatch_value [15:13] : _3541_;
  assign _3545_ = _3846_ ? _0018_[15:13] : 3'h7;
  assign _3547_ = _3834_ ? dscratch1_q[15:13] : dscratch0_q[15:13];
  assign _3549_ = _2017_ ? _3545_ : _3547_;
  assign _3551_ = _0466_ ? _3543_ : _3549_;
  assign _3553_ = _3836_ ? csr_depc_o[15:13] : dcsr_q[15:13];
  assign _3555_ = _3839_ ? mtval_q[15:13] : csr_mepc_o[15:13];
  assign _3557_ = _2011_ ? _3553_ : _3555_;
  assign _3559_ = _3837_ ? csr_mtvec_o[15:13] : mscratch_q[15:13];
  assign _3561_ = _3888_ ? hart_id_i[15:13] : 3'h0;
  assign _3563_ = _1999_ ? _3559_ : _3561_;
  assign _3565_ = _0468_ ? _3557_ : _3563_;
  assign csr_rdata_o[15:13] = _0470_ ? _3551_ : _3565_;
  assign _3567_ = _3742_ ? \gen_trigger_regs.selected_tmatch_value [20:18] : _0016_[52:50];
  assign _3569_ = _3830_ ? _0016_[20:18] : _0018_[20:18];
  assign _3571_ = _1993_ ? _3567_ : _3569_;
  assign _3573_ = _3833_ ? 3'h7 : dscratch1_q[20:18];
  assign _3575_ = _3836_ ? csr_depc_o[20:18] : dcsr_q[20:18];
  assign _3577_ = _3835_ ? dscratch0_q[20:18] : _3575_;
  assign _3579_ = _1995_ ? _3573_ : _3577_;
  assign _3581_ = _0428_ ? _3571_ : _3579_;
  assign _3583_ = _3892_ ? irq_fast_i[4:2] : mtval_q[20:18];
  assign _3585_ = _3841_ ? csr_mepc_o[20:18] : csr_mtvec_o[20:18];
  assign _3587_ = _2003_ ? _3583_ : _3585_;
  assign _3589_ = _3842_ ? mscratch_q[20:18] : mie_q[4:2];
  assign _3591_ = _3888_ ? hart_id_i[20:18] : 3'h0;
  assign _3593_ = _3890_ ? 3'h4 : _3591_;
  assign _3595_ = _2005_ ? _3589_ : _3593_;
  assign _3597_ = _0436_ ? _3587_ : _3595_;
  assign csr_rdata_o[20:18] = _0438_ ? _3581_ : _3597_;
  assign _3599_ = _3742_ ? \gen_trigger_regs.selected_tmatch_value [16] : _0016_[48];
  assign _3601_ = _3830_ ? _0016_[16] : _0018_[16];
  assign _3603_ = _1993_ ? _3599_ : _3601_;
  assign _3605_ = _3833_ ? 1'h1 : dscratch1_q[16];
  assign _3607_ = _3835_ ? dscratch0_q[16] : csr_depc_o[16];
  assign _3609_ = _1995_ ? _3605_ : _3607_;
  assign _3611_ = _0428_ ? _3603_ : _3609_;
  assign _3613_ = _3822_ ? dcsr_q[16] : irq_fast_i[0];
  assign _3615_ = _3839_ ? mtval_q[16] : csr_mepc_o[16];
  assign _3617_ = _2019_ ? _3613_ : _3615_;
  assign _3619_ = _3837_ ? csr_mtvec_o[16] : mscratch_q[16];
  assign _3621_ = _3888_ ? hart_id_i[16] : 1'h0;
  assign _3623_ = _3843_ ? mie_q[0] : _3621_;
  assign _3625_ = _1999_ ? _3619_ : _3623_;
  assign _3627_ = _0472_ ? _3617_ : _3625_;
  assign csr_rdata_o[16] = _0432_ ? _3611_ : _3627_;
  assign _3629_ = _3742_ ? \gen_trigger_regs.selected_tmatch_value [17] : _0016_[49];
  assign _3631_ = _3830_ ? _0016_[17] : _0018_[17];
  assign _3633_ = _1993_ ? _3629_ : _3631_;
  assign _3635_ = _3833_ ? 1'h1 : dscratch1_q[17];
  assign _3637_ = _3836_ ? csr_depc_o[17] : dcsr_q[17];
  assign _3639_ = _3835_ ? dscratch0_q[17] : _3637_;
  assign _3641_ = _1995_ ? _3635_ : _3639_;
  assign _3643_ = _0428_ ? _3633_ : _3641_;
  assign _3645_ = _3892_ ? irq_fast_i[1] : mtval_q[17];
  assign _3647_ = _3841_ ? csr_mepc_o[17] : csr_mtvec_o[17];
  assign _3649_ = _2003_ ? _3645_ : _3647_;
  assign _3651_ = _3842_ ? mscratch_q[17] : mie_q[1];
  assign _3653_ = _3888_ ? hart_id_i[17] : 1'h0;
  assign _3655_ = _3823_ ? mstatus_q[1] : _3653_;
  assign _3657_ = _2005_ ? _3651_ : _3655_;
  assign _3659_ = _0436_ ? _3649_ : _3657_;
  assign csr_rdata_o[17] = _0438_ ? _3643_ : _3659_;
  assign _3661_ = _3832_ ? cpuctrl_q[2:0] : \gen_trigger_regs.selected_tmatch_value [2:0];
  assign _3663_ = _3737_ ? { 2'h0, \gen_trigger_regs.tselect_q  } : _0016_[34:32];
  assign _3665_ = _3740_ ? { \gen_trigger_regs.selected_tmatch_control , 2'h0 } : _3663_;
  assign _3667_ = _2007_ ? _3661_ : _3665_;
  assign _3669_ = _3830_ ? _0016_[2:0] : _0018_[2:0];
  assign _3671_ = _3834_ ? dscratch1_q[2:0] : dscratch0_q[2:0];
  assign _3673_ = _3833_ ? { mcountinhibit[2], 1'h0, mcountinhibit[0] } : _3671_;
  assign _3675_ = _2009_ ? _3669_ : _3673_;
  assign _3677_ = _0474_ ? _3667_ : _3675_;
  assign _3679_ = _3836_ ? csr_depc_o[2:0] : dcsr_q[2:0];
  assign _3681_ = _3840_ ? mcause_q[2:0] : csr_mepc_o[2:0];
  assign _3683_ = _3839_ ? mtval_q[2:0] : _3681_;
  assign _3685_ = _2011_ ? _3679_ : _3683_;
  assign _3687_ = _3837_ ? csr_mtvec_o[2:0] : mscratch_q[2:0];
  assign _3689_ = _3888_ ? hart_id_i[2:0] : 3'h0;
  assign _3691_ = _3890_ ? 3'h4 : _3689_;
  assign _3693_ = _1999_ ? _3687_ : _3691_;
  assign _3695_ = _0476_ ? _3685_ : _3693_;
  assign csr_rdata_o[2:0] = _0478_ ? _3677_ : _3695_;
  assign _3697_ = _3742_ ? \gen_trigger_regs.selected_tmatch_value [12] : 1'h1;
  assign _3699_ = _3826_ ? _0016_[44] : _0016_[12];
  assign _3701_ = _2023_ ? _3697_ : _3699_;
  assign _3703_ = _3846_ ? _0018_[12] : mcountinhibit[12];
  assign _3705_ = _3834_ ? dscratch1_q[12] : dscratch0_q[12];
  assign _3707_ = _2017_ ? _3703_ : _3705_;
  assign _3709_ = _0480_ ? _3701_ : _3707_;
  assign _3711_ = _3836_ ? csr_depc_o[12] : dcsr_q[12];
  assign _3713_ = _3839_ ? mtval_q[12] : csr_mepc_o[12];
  assign _3715_ = _2011_ ? _3711_ : _3713_;
  assign _3717_ = _3837_ ? csr_mtvec_o[12] : mscratch_q[12];
  assign _3719_ = _3888_ ? hart_id_i[12] : 1'h0;
  assign _3721_ = _3823_ ? mstatus_q[3] : _3719_;
  assign _3723_ = _1999_ ? _3717_ : _3721_;
  assign _3725_ = _0468_ ? _3715_ : _3723_;
  assign csr_rdata_o[12] = _0482_ ? _3709_ : _3725_;
  assign _3001_ = _0158_ ? _0371_ : 1'h1;
  assign illegal_csr = _0156_ ? 1'h0 : _3001_;
  assign _0529_ = | _3761_;
  assign _3728_ = $signed(_3760_) < 0 ? 1'h0 << - _3760_ : 1'h0 >> _3760_;
  assign _3762_ = { _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_ } | _3728_;
  assign _3729_ = csr_addr_i[11:10] == 2'h3;
  assign _3739_ = ~ \gen_trigger_regs.tselect_q ;
  assign _3744_ = pc_if_i == \gen_trigger_regs.selected_tmatch_value ;
  assign illegal_csr_priv = csr_addr_i[9:8] > priv_mode_id_o;
  assign illegal_csr_write = _3729_ && csr_wr;
  assign _3746_ = _3752_ && _3754_;
  assign _3748_ = _3756_ && _3758_;
  assign _3750_ = csr_wdata_int < 32'd1;
  assign _3752_ = csr_wdata_int[12:11] != 2'h3;
  assign _3754_ = | csr_wdata_int[12:11];
  assign _3756_ = csr_wdata_int[1:0] != 2'h3;
  assign _3758_ = | csr_wdata_int[1:0];
  assign _3760_ = - $signed({ 27'h0000000, csr_addr_i[4:0] });
  assign _3763_ = ~ illegal_csr_insn_o;
  assign _0121_ = ~ mcountinhibit[0];
  assign _3764_ = ~ mcountinhibit[2];
  assign _3765_ = ~ mcountinhibit[3];
  assign _3766_ = ~ mcountinhibit[4];
  assign _3767_ = ~ mcountinhibit[5];
  assign _3768_ = ~ mcountinhibit[6];
  assign _3769_ = ~ mcountinhibit[7];
  assign _3770_ = ~ mcountinhibit[8];
  assign _3771_ = ~ mcountinhibit[9];
  assign _3772_ = ~ mcountinhibit[10];
  assign _3773_ = ~ mcountinhibit[11];
  assign _3774_ = ~ mcountinhibit[12];
  assign _3063_ = _0115_ | _3966_;
  assign _3776_ = illegal_csr | illegal_csr_write;
  assign _3778_ = _3776_ | illegal_csr_priv;
  assign _3780_ = csr_wdata_i | csr_rdata_o;
  assign _3782_ = mstatus_err | mtvec_err;
  assign csr_shadow_err_o = _3782_ | cpuctrl_err;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) priv_mode_id_o <= 2'h3;
    else priv_mode_id_o <= priv_mode_if_o;
  assign _3784_ = ! csr_op_i;
  assign _3731_ = csr_op_i == 2'h3;
  assign _3733_ = csr_op_i == 2'h2;
  assign _3735_ = csr_op_i == 2'h1;
  assign _3786_ = csr_restore_mret_i ? mstatus_q[4] : _0010_[5];
  assign _3788_ = csr_restore_dret_i ? _0010_[5] : _3786_;
  assign mstatus_d[5] = csr_save_cause_i ? _0097_[3] : _3788_;
  assign _0105_ = nmi_mode_i ? 1'h1 : _0006_;
  assign _0085_ = nmi_mode_i ? mstack_epc_q : { csr_wdata_int[31:1], 1'h0 };
  assign _0107_ = nmi_mode_i ? 1'h1 : _0008_;
  assign _0113_[1:0] = nmi_mode_i ? mstack_q[1:0] : 2'h0;
  assign _0113_[2] = nmi_mode_i ? mstack_q[2] : 1'h1;
  assign _3790_ = csr_restore_mret_i ? _0113_ : _0010_[4:2];
  assign _3792_ = csr_restore_dret_i ? _0010_[4:2] : _3790_;
  assign mstatus_d[4:2] = csr_save_cause_i ? _0097_[2:0] : _3792_;
  assign _0081_ = nmi_mode_i ? mstack_cause_q : { csr_wdata_int[31], csr_wdata_int[4:0] };
  assign _0068_ = debug_mode_i ? { csr_wdata_int[31], csr_wdata_int[4:0] } : csr_mcause_i;
  assign _0093_ = debug_mode_i ? _0006_ : 1'h1;
  assign _0070_ = debug_mode_i ? { csr_wdata_int[31:1], 1'h0 } : _0034_;
  assign _0095_ = debug_mode_i ? _0008_ : 1'h1;
  assign _0072_ = debug_mode_i ? 1'h0 : 1'h1;
  assign _0109_[1:0] = debug_mode_i ? _0010_[3:2] : priv_mode_id_o;
  assign _0109_[2] = debug_mode_i ? _0010_[4] : mstatus_q[5];
  assign _0099_ = debug_mode_i ? _0012_ : 1'h1;
  assign _0075_ = debug_mode_i ? csr_wdata_int : csr_mtval_i;
  assign _0101_ = debug_mode_i ? _0014_ : 1'h1;
  assign _0079_ = debug_csr_save_i ? 1'h1 : _0004_;
  assign _0026_ = debug_csr_save_i ? _0034_ : { csr_wdata_int[31:1], 1'h0 };
  assign _0077_ = debug_csr_save_i ? 1'h1 : _0002_;
  assign _0111_ = debug_csr_save_i ? debug_cause_i : _0000_[8:6];
  assign _0103_ = debug_csr_save_i ? priv_mode_id_o : _0000_[1:0];
  assign _0054_ = debug_csr_save_i ? 1'h0 : _0072_;
  assign _0091_ = debug_csr_save_i ? _0014_ : _0101_;
  assign _0060_ = debug_csr_save_i ? csr_wdata_int : _0075_;
  assign _0083_ = debug_csr_save_i ? _0006_ : _0093_;
  assign _0036_ = debug_csr_save_i ? { csr_wdata_int[31], csr_wdata_int[4:0] } : _0068_;
  assign _0087_ = debug_csr_save_i ? _0008_ : _0095_;
  assign _0042_ = debug_csr_save_i ? { csr_wdata_int[31:1], 1'h0 } : _0070_;
  assign _0089_ = debug_csr_save_i ? _0012_ : _0099_;
  assign _0097_ = debug_csr_save_i ? _0010_[5:2] : _0109_;
  assign _3794_ = csr_save_wb_i ? pc_wb_i : pc_id_i;
  assign _3796_ = csr_save_id_i ? pc_id_i : _3794_;
  assign _0034_ = csr_save_if_i ? pc_if_i : _3796_;
  assign mstack_en = csr_save_cause_i ? _0054_ : 1'h0;
  assign depc_en = csr_save_cause_i ? _0079_ : _0004_;
  assign depc_d = csr_save_cause_i ? _0026_ : { csr_wdata_int[31:1], 1'h0 };
  assign dcsr_en = csr_save_cause_i ? _0077_ : _0002_;
  assign dcsr_d[8:6] = csr_save_cause_i ? _0111_ : _0000_[8:6];
  assign dcsr_d[1:0] = csr_save_cause_i ? _0103_ : _0000_[1:0];
  assign mtval_en = csr_save_cause_i ? _0091_ : _0014_;
  assign mtval_d = csr_save_cause_i ? _0060_ : csr_wdata_int;
  assign _3798_ = csr_restore_mret_i ? _0105_ : _0006_;
  assign _3800_ = csr_restore_dret_i ? _0006_ : _3798_;
  assign mcause_en = csr_save_cause_i ? _0083_ : _3800_;
  assign _3802_ = csr_restore_mret_i ? _0081_ : { csr_wdata_int[31], csr_wdata_int[4:0] };
  assign _3804_ = csr_restore_dret_i ? { csr_wdata_int[31], csr_wdata_int[4:0] } : _3802_;
  assign mcause_d = csr_save_cause_i ? _0036_ : _3804_;
  assign _3806_ = csr_restore_mret_i ? _0107_ : _0008_;
  assign _3808_ = csr_restore_dret_i ? _0008_ : _3806_;
  assign mepc_en = csr_save_cause_i ? _0087_ : _3808_;
  assign _3810_ = csr_restore_mret_i ? _0085_ : { csr_wdata_int[31:1], 1'h0 };
  assign _3812_ = csr_restore_dret_i ? { csr_wdata_int[31:1], 1'h0 } : _3810_;
  assign mepc_d = csr_save_cause_i ? _0042_ : _3812_;
  assign _3814_ = csr_restore_mret_i ? 1'h1 : _0012_;
  assign _3816_ = csr_restore_dret_i ? _0012_ : _3814_;
  assign mstatus_en = csr_save_cause_i ? _0089_ : _3816_;
  assign _0109_[3] = debug_mode_i ? _0010_[5] : 1'h0;
  assign _3818_ = csr_restore_mret_i ? mstatus_q[3:2] : priv_mode_id_o;
  assign _3820_ = csr_restore_dret_i ? dcsr_q[1:0] : _3818_;
  assign priv_mode_if_o = csr_save_cause_i ? 2'h3 : _3820_;
  assign _0022_[31:28] = _3822_ ? 4'h4 : dcsr_q[31:28];
  assign _0056_[5:4] = _3823_ ? { csr_wdata_int[3], csr_wdata_int[7] } : mstatus_q[5:4];
  assign _0056_[3:2] = _3823_ ? _0073_ : mstatus_q[3:2];
  assign _0022_[15] = _3822_ ? csr_wdata_int[15] : dcsr_q[15];
  assign _0022_[14] = _3822_ ? 1'h0 : dcsr_q[14];
  assign _0022_[27:16] = _3822_ ? 12'h000 : dcsr_q[27:16];
  assign _0056_[1:0] = _3823_ ? { csr_wdata_int[17], csr_wdata_int[21] } : mstatus_q[1:0];
  assign _0022_[1:0] = _3822_ ? _0066_ : dcsr_q[1:0];
  assign _0022_[5] = _3822_ ? 1'h0 : dcsr_q[5];
  assign _0022_[4] = _3822_ ? 1'h0 : dcsr_q[4];
  assign _0022_[3] = _3822_ ? 1'h0 : dcsr_q[3];
  assign _0022_[2] = _3822_ ? csr_wdata_int[2] : dcsr_q[2];
  assign _0022_[13:12] = _3822_ ? csr_wdata_int[13:12] : dcsr_q[13:12];
  assign _0022_[11] = _3822_ ? 1'h0 : dcsr_q[11];
  assign _0066_ = _3748_ ? 2'h3 : csr_wdata_int[1:0];
  assign _0022_[9] = _3822_ ? 1'h0 : dcsr_q[9];
  assign _0073_ = _3746_ ? 2'h3 : csr_wdata_int[12:11];
  assign _0058_ = _3823_ ? 1'h1 : 1'h0;
  assign _0020_ = _3832_ ? 1'h1 : 1'h0;
  assign _0048_ = _3826_ ? _3063_ : 32'd0;
  assign _0046_ = _3830_ ? _3063_ : 32'd0;
  assign _0040_ = _3833_ ? 1'h1 : 1'h0;
  assign _0032_ = _3834_ ? 1'h1 : 1'h0;
  assign _0030_ = _3835_ ? 1'h1 : 1'h0;
  assign _0028_ = _3836_ ? 1'h1 : 1'h0;
  assign _0024_ = _3822_ ? 1'h1 : 1'h0;
  assign _0022_[10] = _3822_ ? 1'h0 : dcsr_q[10];
  assign _0064_ = _3837_ ? 1'h1 : csr_mtvec_init_i;
  assign _0062_ = _3839_ ? 1'h1 : 1'h0;
  assign _0038_ = _3840_ ? 1'h1 : 1'h0;
  assign _0044_ = _3841_ ? 1'h1 : 1'h0;
  assign _0052_ = _3842_ ? 1'h1 : 1'h0;
  assign _0050_ = _3843_ ? 1'h1 : 1'h0;
  assign cpuctrl_we = csr_we_int ? _0020_ : 1'h0;
  assign mhpmcounterh_we = csr_we_int ? _0048_ : 32'd0;
  assign mhpmcounter_we = csr_we_int ? _0046_ : 32'd0;
  assign mcountinhibit_we = csr_we_int ? _0040_ : 1'h0;
  assign dscratch1_en = csr_we_int ? _0032_ : 1'h0;
  assign dscratch0_en = csr_we_int ? _0030_ : 1'h0;
  assign _0004_ = csr_we_int ? _0028_ : 1'h0;
  assign _0002_ = csr_we_int ? _0024_ : 1'h0;
  assign { dcsr_d[31:9], _0000_[8:6], dcsr_d[5:2], _0000_[1:0] } = csr_we_int ? { _0022_[31:9], dcsr_q[8:6], _0022_[5:0] } : dcsr_q;
  assign mtvec_en = csr_we_int ? _0064_ : csr_mtvec_init_i;
  assign _0014_ = csr_we_int ? _0062_ : 1'h0;
  assign _0006_ = csr_we_int ? _0038_ : 1'h0;
  assign _0008_ = csr_we_int ? _0044_ : 1'h0;
  assign mscratch_en = csr_we_int ? _0052_ : 1'h0;
  assign mie_en = csr_we_int ? _0050_ : 1'h0;
  assign _0012_ = csr_we_int ? _0058_ : 1'h0;
  assign { _0010_[5:2], mstatus_d[1:0] } = csr_we_int ? _0056_ : mstatus_q;
  assign _3826_ = | _3824_;
  assign _3846_ = | _3844_;
  assign _3892_ = csr_addr_i == 12'h344;
  assign _3843_ = csr_addr_i == 12'h304;
  assign _3894_ = csr_addr_i[4:0] == 5'h1f;
  assign _3896_ = csr_addr_i[4:0] == 5'h1e;
  assign _3898_ = csr_addr_i[4:0] == 5'h1d;
  assign _3900_ = csr_addr_i[4:0] == 5'h1c;
  assign _3902_ = csr_addr_i[4:0] == 5'h1b;
  assign _3904_ = csr_addr_i[4:0] == 5'h1a;
  assign _3906_ = csr_addr_i[4:0] == 5'h19;
  assign _3908_ = csr_addr_i[4:0] == 5'h18;
  assign _3910_ = csr_addr_i[4:0] == 5'h17;
  assign _3912_ = csr_addr_i[4:0] == 5'h16;
  assign _3914_ = csr_addr_i[4:0] == 5'h15;
  assign _3916_ = csr_addr_i[4:0] == 5'h14;
  assign _3918_ = csr_addr_i[4:0] == 5'h13;
  assign _3920_ = csr_addr_i[4:0] == 5'h12;
  assign _3922_ = csr_addr_i[4:0] == 5'h11;
  assign _3924_ = csr_addr_i[4:0] == 5'h10;
  assign _3926_ = csr_addr_i[4:0] == 5'h0f;
  assign _3928_ = csr_addr_i[4:0] == 5'h0e;
  assign _3930_ = csr_addr_i[4:0] == 5'h0d;
  assign _3932_ = csr_addr_i[4:0] == 5'h0c;
  assign _3934_ = csr_addr_i[4:0] == 5'h0b;
  assign _3936_ = csr_addr_i[4:0] == 5'h0a;
  assign _3938_ = csr_addr_i[4:0] == 5'h09;
  assign _3940_ = csr_addr_i[4:0] == 5'h08;
  assign _3942_ = csr_addr_i[4:0] == 5'h07;
  assign _3944_ = csr_addr_i[4:0] == 5'h06;
  assign _3946_ = csr_addr_i[4:0] == 5'h05;
  assign _3948_ = csr_addr_i[4:0] == 5'h04;
  assign _3950_ = csr_addr_i[4:0] == 5'h03;
  assign _3952_ = csr_addr_i[4:0] == 5'h02;
  assign _3954_ = csr_addr_i[4:0] == 5'h01;
  assign _3840_ = csr_addr_i == 12'h342;
  assign _3833_ = csr_addr_i == 12'h320;
  assign _3834_ = csr_addr_i == 12'h7b3;
  assign _3835_ = csr_addr_i == 12'h7b2;
  assign _3836_ = csr_addr_i == 12'h7b1;
  assign _3822_ = csr_addr_i == 12'h7b0;
  assign _3848_ = csr_addr_i == 12'h3bf;
  assign _3850_ = csr_addr_i == 12'h3be;
  assign _3852_ = csr_addr_i == 12'h3bd;
  assign _3854_ = csr_addr_i == 12'h3bc;
  assign _3856_ = csr_addr_i == 12'h3bb;
  assign _3858_ = csr_addr_i == 12'h3ba;
  assign _3860_ = csr_addr_i == 12'h3b9;
  assign _3862_ = csr_addr_i == 12'h3b8;
  assign _3864_ = csr_addr_i == 12'h3b7;
  assign _3866_ = csr_addr_i == 12'h3b6;
  assign _3868_ = csr_addr_i == 12'h3b5;
  assign _3870_ = csr_addr_i == 12'h3b4;
  assign _3872_ = csr_addr_i == 12'h3b3;
  assign _3874_ = csr_addr_i == 12'h3b2;
  assign _3876_ = csr_addr_i == 12'h3b1;
  assign _3878_ = csr_addr_i == 12'h3b0;
  assign _3880_ = csr_addr_i == 12'h3a3;
  assign _3882_ = csr_addr_i == 12'h3a2;
  assign _3884_ = csr_addr_i == 12'h3a1;
  assign _3886_ = csr_addr_i == 12'h3a0;
  assign _3839_ = csr_addr_i == 12'h343;
  assign _3841_ = csr_addr_i == 12'h341;
  assign _3837_ = csr_addr_i == 12'h305;
  assign _3842_ = csr_addr_i == 12'h340;
  assign _3890_ = csr_addr_i == 12'h301;
  assign _3823_ = csr_addr_i == 12'h300;
  assign _3888_ = csr_addr_i == 12'hf14;
  assign _3830_ = | _3828_;
  assign _3828_[18] = csr_addr_i == 12'hb13;
  assign _3828_[19] = csr_addr_i == 12'hb14;
  assign _3828_[20] = csr_addr_i == 12'hb15;
  assign _3828_[21] = csr_addr_i == 12'hb16;
  assign _3828_[22] = csr_addr_i == 12'hb17;
  assign _3828_[23] = csr_addr_i == 12'hb18;
  assign _3828_[24] = csr_addr_i == 12'hb19;
  assign _3828_[25] = csr_addr_i == 12'hb1a;
  assign _3828_[26] = csr_addr_i == 12'hb1b;
  assign _3828_[27] = csr_addr_i == 12'hb1c;
  assign _3828_[28] = csr_addr_i == 12'hb1d;
  assign _3828_[29] = csr_addr_i == 12'hb1e;
  assign _3828_[30] = csr_addr_i == 12'hb1f;
  assign _3844_[0] = csr_addr_i == 12'h323;
  assign _3844_[1] = csr_addr_i == 12'h324;
  assign _3844_[10] = csr_addr_i == 12'h32d;
  assign _3844_[11] = csr_addr_i == 12'h32e;
  assign _3844_[12] = csr_addr_i == 12'h32f;
  assign _3844_[13] = csr_addr_i == 12'h330;
  assign _3844_[14] = csr_addr_i == 12'h331;
  assign _3844_[15] = csr_addr_i == 12'h332;
  assign _3844_[16] = csr_addr_i == 12'h333;
  assign _3844_[17] = csr_addr_i == 12'h334;
  assign _3844_[18] = csr_addr_i == 12'h335;
  assign _3844_[19] = csr_addr_i == 12'h336;
  assign _3844_[2] = csr_addr_i == 12'h325;
  assign _3844_[20] = csr_addr_i == 12'h337;
  assign _3844_[21] = csr_addr_i == 12'h338;
  assign _3844_[22] = csr_addr_i == 12'h339;
  assign _3844_[23] = csr_addr_i == 12'h33a;
  assign _3844_[24] = csr_addr_i == 12'h33b;
  assign _3844_[25] = csr_addr_i == 12'h33c;
  assign _3844_[26] = csr_addr_i == 12'h33d;
  assign _3844_[27] = csr_addr_i == 12'h33e;
  assign _3844_[28] = csr_addr_i == 12'h33f;
  assign _3844_[3] = csr_addr_i == 12'h326;
  assign _3844_[4] = csr_addr_i == 12'h327;
  assign _3844_[5] = csr_addr_i == 12'h328;
  assign _3844_[6] = csr_addr_i == 12'h329;
  assign _3844_[7] = csr_addr_i == 12'h32a;
  assign _3844_[8] = csr_addr_i == 12'h32b;
  assign _3844_[9] = csr_addr_i == 12'h32c;
  assign _3956_ = csr_addr_i == 12'h7c1;
  assign _3832_ = csr_addr_i == 12'h7c0;
  assign _3958_ = csr_addr_i == 12'h7aa;
  assign _3960_ = csr_addr_i == 12'h7a8;
  assign _3962_ = csr_addr_i == 12'h7a3;
  assign _3742_ = csr_addr_i == 12'h7a2;
  assign _3740_ = csr_addr_i == 12'h7a1;
  assign _3737_ = csr_addr_i == 12'h7a0;
  assign _3824_[0] = csr_addr_i == 12'hb80;
  assign _3824_[1] = csr_addr_i == 12'hb82;
  assign _3824_[10] = csr_addr_i == 12'hb8b;
  assign _3824_[11] = csr_addr_i == 12'hb8c;
  assign _3824_[12] = csr_addr_i == 12'hb8d;
  assign _3824_[13] = csr_addr_i == 12'hb8e;
  assign _3824_[14] = csr_addr_i == 12'hb8f;
  assign _3824_[15] = csr_addr_i == 12'hb90;
  assign _3824_[16] = csr_addr_i == 12'hb91;
  assign _3824_[17] = csr_addr_i == 12'hb92;
  assign _3824_[18] = csr_addr_i == 12'hb93;
  assign _3824_[19] = csr_addr_i == 12'hb94;
  assign _3824_[2] = csr_addr_i == 12'hb83;
  assign _3824_[20] = csr_addr_i == 12'hb95;
  assign _3824_[21] = csr_addr_i == 12'hb96;
  assign _3824_[22] = csr_addr_i == 12'hb97;
  assign _3824_[23] = csr_addr_i == 12'hb98;
  assign _3824_[24] = csr_addr_i == 12'hb99;
  assign _3824_[25] = csr_addr_i == 12'hb9a;
  assign _3824_[26] = csr_addr_i == 12'hb9b;
  assign _3824_[27] = csr_addr_i == 12'hb9c;
  assign _3824_[28] = csr_addr_i == 12'hb9d;
  assign _3824_[29] = csr_addr_i == 12'hb9e;
  assign _3824_[3] = csr_addr_i == 12'hb84;
  assign _3824_[30] = csr_addr_i == 12'hb9f;
  assign _3824_[4] = csr_addr_i == 12'hb85;
  assign _3824_[5] = csr_addr_i == 12'hb86;
  assign _3824_[6] = csr_addr_i == 12'hb87;
  assign _3824_[7] = csr_addr_i == 12'hb88;
  assign _3824_[8] = csr_addr_i == 12'hb89;
  assign _3824_[9] = csr_addr_i == 12'hb8a;
  assign _3828_[0] = csr_addr_i == 12'hb00;
  assign _3828_[1] = csr_addr_i == 12'hb02;
  assign _3828_[10] = csr_addr_i == 12'hb0b;
  assign _3828_[11] = csr_addr_i == 12'hb0c;
  assign _3828_[12] = csr_addr_i == 12'hb0d;
  assign _3828_[13] = csr_addr_i == 12'hb0e;
  assign _3828_[14] = csr_addr_i == 12'hb0f;
  assign _3828_[15] = csr_addr_i == 12'hb10;
  assign _3828_[16] = csr_addr_i == 12'hb11;
  assign _3828_[17] = csr_addr_i == 12'hb12;
  assign _3828_[2] = csr_addr_i == 12'hb03;
  assign _3828_[3] = csr_addr_i == 12'hb04;
  assign _3828_[4] = csr_addr_i == 12'hb05;
  assign _3828_[5] = csr_addr_i == 12'hb06;
  assign _3828_[6] = csr_addr_i == 12'hb07;
  assign _3828_[7] = csr_addr_i == 12'hb08;
  assign _3828_[8] = csr_addr_i == 12'hb09;
  assign _3828_[9] = csr_addr_i == 12'hb0a;
  assign _3964_ = csr_addr_i == 12'h306;
  assign csr_wr = | { _3735_, _3733_, _3731_ };
  assign irq_pending_o = | irqs_o;
  assign _3966_ = $signed(_3760_) < 0 ? 1'h1 << - _3760_ : 1'h1 >> _3760_;
  assign mtvec_d = csr_mtvec_init_i ? { boot_addr_i[31:8], 8'h01 } : { csr_wdata_int[31:8], 8'h01 };
  assign priv_mode_lsu_o = mstatus_q[1] ? mstatus_q[3:2] : priv_mode_id_o;
  assign \gen_trigger_regs.tselect_d  = _3750_ ? csr_wdata_int[0] : 1'h0;
  paramodauxy_ibex_counterCounterWidth3200000000000000000000000000100000  \gen_cntrs[0].gen_imp.mcounters_variable_i  (
    .clk_i(clk_i),
    .counter_inc_i(_0124_),
    .counter_inc_i_t0(_0125_),
    .counter_val_i(csr_wdata_int),
    .counter_val_i_t0(csr_wdata_int_t0),
    .counter_val_o(\mhpmcounter[3] ),
    .counter_val_o_t0(\mhpmcounter[3]_t0 ),
    .counter_we_i(mhpmcounter_we[3]),
    .counter_we_i_t0(mhpmcounter_we_t0[3]),
    .counterh_we_i(mhpmcounterh_we[3]),
    .counterh_we_i_t0(mhpmcounterh_we_t0[3]),
    .rst_ni(rst_ni)
  );
  paramodauxy_ibex_counterCounterWidth3200000000000000000000000000100000  \gen_cntrs[1].gen_imp.mcounters_variable_i  (
    .clk_i(clk_i),
    .counter_inc_i(_0126_),
    .counter_inc_i_t0(_0127_),
    .counter_val_i(csr_wdata_int),
    .counter_val_i_t0(csr_wdata_int_t0),
    .counter_val_o(\mhpmcounter[4] ),
    .counter_val_o_t0(\mhpmcounter[4]_t0 ),
    .counter_we_i(mhpmcounter_we[4]),
    .counter_we_i_t0(mhpmcounter_we_t0[4]),
    .counterh_we_i(mhpmcounterh_we[4]),
    .counterh_we_i_t0(mhpmcounterh_we_t0[4]),
    .rst_ni(rst_ni)
  );
  paramodauxy_ibex_counterCounterWidth3200000000000000000000000000100000  \gen_cntrs[2].gen_imp.mcounters_variable_i  (
    .clk_i(clk_i),
    .counter_inc_i(_0128_),
    .counter_inc_i_t0(_0129_),
    .counter_val_i(csr_wdata_int),
    .counter_val_i_t0(csr_wdata_int_t0),
    .counter_val_o(\mhpmcounter[5] ),
    .counter_val_o_t0(\mhpmcounter[5]_t0 ),
    .counter_we_i(mhpmcounter_we[5]),
    .counter_we_i_t0(mhpmcounter_we_t0[5]),
    .counterh_we_i(mhpmcounterh_we[5]),
    .counterh_we_i_t0(mhpmcounterh_we_t0[5]),
    .rst_ni(rst_ni)
  );
  paramodauxy_ibex_counterCounterWidth3200000000000000000000000000100000  \gen_cntrs[3].gen_imp.mcounters_variable_i  (
    .clk_i(clk_i),
    .counter_inc_i(_0130_),
    .counter_inc_i_t0(_0131_),
    .counter_val_i(csr_wdata_int),
    .counter_val_i_t0(csr_wdata_int_t0),
    .counter_val_o(\mhpmcounter[6] ),
    .counter_val_o_t0(\mhpmcounter[6]_t0 ),
    .counter_we_i(mhpmcounter_we[6]),
    .counter_we_i_t0(mhpmcounter_we_t0[6]),
    .counterh_we_i(mhpmcounterh_we[6]),
    .counterh_we_i_t0(mhpmcounterh_we_t0[6]),
    .rst_ni(rst_ni)
  );
  paramodauxy_ibex_counterCounterWidth3200000000000000000000000000100000  \gen_cntrs[4].gen_imp.mcounters_variable_i  (
    .clk_i(clk_i),
    .counter_inc_i(_0132_),
    .counter_inc_i_t0(_0133_),
    .counter_val_i(csr_wdata_int),
    .counter_val_i_t0(csr_wdata_int_t0),
    .counter_val_o(\mhpmcounter[7] ),
    .counter_val_o_t0(\mhpmcounter[7]_t0 ),
    .counter_we_i(mhpmcounter_we[7]),
    .counter_we_i_t0(mhpmcounter_we_t0[7]),
    .counterh_we_i(mhpmcounterh_we[7]),
    .counterh_we_i_t0(mhpmcounterh_we_t0[7]),
    .rst_ni(rst_ni)
  );
  paramodauxy_ibex_counterCounterWidth3200000000000000000000000000100000  \gen_cntrs[5].gen_imp.mcounters_variable_i  (
    .clk_i(clk_i),
    .counter_inc_i(_0134_),
    .counter_inc_i_t0(_0135_),
    .counter_val_i(csr_wdata_int),
    .counter_val_i_t0(csr_wdata_int_t0),
    .counter_val_o(\mhpmcounter[8] ),
    .counter_val_o_t0(\mhpmcounter[8]_t0 ),
    .counter_we_i(mhpmcounter_we[8]),
    .counter_we_i_t0(mhpmcounter_we_t0[8]),
    .counterh_we_i(mhpmcounterh_we[8]),
    .counterh_we_i_t0(mhpmcounterh_we_t0[8]),
    .rst_ni(rst_ni)
  );
  paramodauxy_ibex_counterCounterWidth3200000000000000000000000000100000  \gen_cntrs[6].gen_imp.mcounters_variable_i  (
    .clk_i(clk_i),
    .counter_inc_i(_0136_),
    .counter_inc_i_t0(_0137_),
    .counter_val_i(csr_wdata_int),
    .counter_val_i_t0(csr_wdata_int_t0),
    .counter_val_o(\mhpmcounter[9] ),
    .counter_val_o_t0(\mhpmcounter[9]_t0 ),
    .counter_we_i(mhpmcounter_we[9]),
    .counter_we_i_t0(mhpmcounter_we_t0[9]),
    .counterh_we_i(mhpmcounterh_we[9]),
    .counterh_we_i_t0(mhpmcounterh_we_t0[9]),
    .rst_ni(rst_ni)
  );
  paramodauxy_ibex_counterCounterWidth3200000000000000000000000000100000  \gen_cntrs[7].gen_imp.mcounters_variable_i  (
    .clk_i(clk_i),
    .counter_inc_i(_0138_),
    .counter_inc_i_t0(_0139_),
    .counter_val_i(csr_wdata_int),
    .counter_val_i_t0(csr_wdata_int_t0),
    .counter_val_o(\mhpmcounter[10] ),
    .counter_val_o_t0(\mhpmcounter[10]_t0 ),
    .counter_we_i(mhpmcounter_we[10]),
    .counter_we_i_t0(mhpmcounter_we_t0[10]),
    .counterh_we_i(mhpmcounterh_we[10]),
    .counterh_we_i_t0(mhpmcounterh_we_t0[10]),
    .rst_ni(rst_ni)
  );
  paramodauxy_ibex_counterCounterWidth3200000000000000000000000000100000  \gen_cntrs[8].gen_imp.mcounters_variable_i  (
    .clk_i(clk_i),
    .counter_inc_i(_0140_),
    .counter_inc_i_t0(_0141_),
    .counter_val_i(csr_wdata_int),
    .counter_val_i_t0(csr_wdata_int_t0),
    .counter_val_o(\mhpmcounter[11] ),
    .counter_val_o_t0(\mhpmcounter[11]_t0 ),
    .counter_we_i(mhpmcounter_we[11]),
    .counter_we_i_t0(mhpmcounter_we_t0[11]),
    .counterh_we_i(mhpmcounterh_we[11]),
    .counterh_we_i_t0(mhpmcounterh_we_t0[11]),
    .rst_ni(rst_ni)
  );
  paramodauxy_ibex_counterCounterWidth3200000000000000000000000000100000  \gen_cntrs[9].gen_imp.mcounters_variable_i  (
    .clk_i(clk_i),
    .counter_inc_i(_0142_),
    .counter_inc_i_t0(_0143_),
    .counter_val_i(csr_wdata_int),
    .counter_val_i_t0(csr_wdata_int_t0),
    .counter_val_o(\mhpmcounter[12] ),
    .counter_val_o_t0(\mhpmcounter[12]_t0 ),
    .counter_we_i(mhpmcounter_we[12]),
    .counter_we_i_t0(mhpmcounter_we_t0[12]),
    .counterh_we_i(mhpmcounterh_we[12]),
    .counterh_we_i_t0(mhpmcounterh_we_t0[12]),
    .rst_ni(rst_ni)
  );
  paramodbc034ef4e1b4bac0b496e4b04aec5350c1a23f8cauxy_ibex_csr  \gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_control_csr  (
    .clk_i(clk_i),
    .rd_data_o(\gen_trigger_regs.selected_tmatch_control ),
    .rd_data_o_t0(\gen_trigger_regs.selected_tmatch_control_t0 ),
    .rst_ni(rst_ni),
    .wr_data_i(csr_wdata_int[2]),
    .wr_data_i_t0(csr_wdata_int_t0[2]),
    .wr_en_i(\gen_trigger_regs.tmatch_control_we ),
    .wr_en_i_t0(\gen_trigger_regs.tmatch_control_we_t0 )
  );
  paramod85ba01ab5a28334786aba5877c1fe04472f39fbaauxy_ibex_csr  \gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr  (
    .clk_i(clk_i),
    .rd_data_o(\gen_trigger_regs.selected_tmatch_value ),
    .rd_data_o_t0(\gen_trigger_regs.selected_tmatch_value_t0 ),
    .rst_ni(rst_ni),
    .wr_data_i(csr_wdata_int),
    .wr_data_i_t0(csr_wdata_int_t0),
    .wr_en_i(\gen_trigger_regs.tmatch_value_we ),
    .wr_en_i_t0(\gen_trigger_regs.tmatch_value_we_t0 )
  );
  paramodeccb28a0d9c7c379466a9299a8885e9ec9033585auxy_ibex_csr  \gen_trigger_regs.u_tselect_csr  (
    .clk_i(clk_i),
    .rd_data_o(\gen_trigger_regs.tselect_q ),
    .rd_data_o_t0(\gen_trigger_regs.tselect_q_t0 ),
    .rst_ni(rst_ni),
    .wr_data_i(\gen_trigger_regs.tselect_d ),
    .wr_data_i_t0(\gen_trigger_regs.tselect_d_t0 ),
    .wr_en_i(\gen_trigger_regs.tselect_we ),
    .wr_en_i_t0(\gen_trigger_regs.tselect_we_t0 )
  );
  paramodauxy_ibex_counterCounterWidths3200000000000000000000000001000000  mcycle_counter_i (
    .clk_i(clk_i),
    .counter_inc_i(_0121_),
    .counter_inc_i_t0(mcountinhibit_t0[0]),
    .counter_val_i(csr_wdata_int),
    .counter_val_i_t0(csr_wdata_int_t0),
    .counter_val_o(\mhpmcounter[0] ),
    .counter_val_o_t0(\mhpmcounter[0]_t0 ),
    .counter_we_i(mhpmcounter_we[0]),
    .counter_we_i_t0(mhpmcounter_we_t0[0]),
    .counterh_we_i(mhpmcounterh_we[0]),
    .counterh_we_i_t0(mhpmcounterh_we_t0[0]),
    .rst_ni(rst_ni)
  );
  paramodauxy_ibex_counterCounterWidths3200000000000000000000000001000000  minstret_counter_i (
    .clk_i(clk_i),
    .counter_inc_i(_0122_),
    .counter_inc_i_t0(_0123_),
    .counter_val_i(csr_wdata_int),
    .counter_val_i_t0(csr_wdata_int_t0),
    .counter_val_o(\mhpmcounter[2] ),
    .counter_val_o_t0(\mhpmcounter[2]_t0 ),
    .counter_we_i(mhpmcounter_we[2]),
    .counter_we_i_t0(mhpmcounter_we_t0[2]),
    .counterh_we_i(mhpmcounterh_we[2]),
    .counterh_we_i_t0(mhpmcounterh_we_t0[2]),
    .rst_ni(rst_ni)
  );
  paramod2736aa8a03348385795fda019fbdaaafd7f2ecf9auxy_ibex_csr  u_cpuctrl_csr (
    .clk_i(clk_i),
    .rd_data_o(cpuctrl_q),
    .rd_data_o_t0(cpuctrl_q_t0),
    .rd_error_o(cpuctrl_err),
    .rd_error_o_t0(cpuctrl_err_t0),
    .rst_ni(rst_ni),
    .wr_data_i(6'h00),
    .wr_data_i_t0(6'h00),
    .wr_en_i(cpuctrl_we),
    .wr_en_i_t0(cpuctrl_we_t0)
  );
  paramod9a435d8f6db004a67362aa9a56f32ea481a74dbeauxy_ibex_csr  u_dcsr_csr (
    .clk_i(clk_i),
    .rd_data_o(dcsr_q),
    .rd_data_o_t0(dcsr_q_t0),
    .rst_ni(rst_ni),
    .wr_data_i(dcsr_d),
    .wr_data_i_t0(dcsr_d_t0),
    .wr_en_i(dcsr_en),
    .wr_en_i_t0(dcsr_en_t0)
  );
  paramod85ba01ab5a28334786aba5877c1fe04472f39fbaauxy_ibex_csr  u_depc_csr (
    .clk_i(clk_i),
    .rd_data_o(csr_depc_o),
    .rd_data_o_t0(csr_depc_o_t0),
    .rst_ni(rst_ni),
    .wr_data_i(depc_d),
    .wr_data_i_t0(depc_d_t0),
    .wr_en_i(depc_en),
    .wr_en_i_t0(depc_en_t0)
  );
  paramod85ba01ab5a28334786aba5877c1fe04472f39fbaauxy_ibex_csr  u_dscratch0_csr (
    .clk_i(clk_i),
    .rd_data_o(dscratch0_q),
    .rd_data_o_t0(dscratch0_q_t0),
    .rst_ni(rst_ni),
    .wr_data_i(csr_wdata_int),
    .wr_data_i_t0(csr_wdata_int_t0),
    .wr_en_i(dscratch0_en),
    .wr_en_i_t0(dscratch0_en_t0)
  );
  paramod85ba01ab5a28334786aba5877c1fe04472f39fbaauxy_ibex_csr  u_dscratch1_csr (
    .clk_i(clk_i),
    .rd_data_o(dscratch1_q),
    .rd_data_o_t0(dscratch1_q_t0),
    .rst_ni(rst_ni),
    .wr_data_i(csr_wdata_int),
    .wr_data_i_t0(csr_wdata_int_t0),
    .wr_en_i(dscratch1_en),
    .wr_en_i_t0(dscratch1_en_t0)
  );
  paramod2736aa8a03348385795fda019fbdaaafd7f2ecf9auxy_ibex_csr  u_mcause_csr (
    .clk_i(clk_i),
    .rd_data_o(mcause_q),
    .rd_data_o_t0(mcause_q_t0),
    .rst_ni(rst_ni),
    .wr_data_i(mcause_d),
    .wr_data_i_t0(mcause_d_t0),
    .wr_en_i(mcause_en),
    .wr_en_i_t0(mcause_en_t0)
  );
  paramod85ba01ab5a28334786aba5877c1fe04472f39fbaauxy_ibex_csr  u_mepc_csr (
    .clk_i(clk_i),
    .rd_data_o(csr_mepc_o),
    .rd_data_o_t0(csr_mepc_o_t0),
    .rst_ni(rst_ni),
    .wr_data_i(mepc_d),
    .wr_data_i_t0(mepc_d_t0),
    .wr_en_i(mepc_en),
    .wr_en_i_t0(mepc_en_t0)
  );
  paramode55993a14b1fbc43320d549f521b710ed37596c6auxy_ibex_csr  u_mie_csr (
    .clk_i(clk_i),
    .rd_data_o(mie_q),
    .rd_data_o_t0(mie_q_t0),
    .rst_ni(rst_ni),
    .wr_data_i({ csr_wdata_int[3], csr_wdata_int[7], csr_wdata_int[11], csr_wdata_int[30:16] }),
    .wr_data_i_t0({ csr_wdata_int_t0[3], csr_wdata_int_t0[7], csr_wdata_int_t0[11], csr_wdata_int_t0[30:16] }),
    .wr_en_i(mie_en),
    .wr_en_i_t0(mie_en_t0)
  );
  paramod85ba01ab5a28334786aba5877c1fe04472f39fbaauxy_ibex_csr  u_mscratch_csr (
    .clk_i(clk_i),
    .rd_data_o(mscratch_q),
    .rd_data_o_t0(mscratch_q_t0),
    .rst_ni(rst_ni),
    .wr_data_i(csr_wdata_int),
    .wr_data_i_t0(csr_wdata_int_t0),
    .wr_en_i(mscratch_en),
    .wr_en_i_t0(mscratch_en_t0)
  );
  paramod2736aa8a03348385795fda019fbdaaafd7f2ecf9auxy_ibex_csr  u_mstack_cause_csr (
    .clk_i(clk_i),
    .rd_data_o(mstack_cause_q),
    .rd_data_o_t0(mstack_cause_q_t0),
    .rst_ni(rst_ni),
    .wr_data_i(mcause_q),
    .wr_data_i_t0(mcause_q_t0),
    .wr_en_i(mstack_en),
    .wr_en_i_t0(mstack_en_t0)
  );
  paramod410b37fbfbfa994790f1902c150d2be939cadb3bauxy_ibex_csr  u_mstack_csr (
    .clk_i(clk_i),
    .rd_data_o(mstack_q),
    .rd_data_o_t0(mstack_q_t0),
    .rst_ni(rst_ni),
    .wr_data_i(mstatus_q[4:2]),
    .wr_data_i_t0(mstatus_q_t0[4:2]),
    .wr_en_i(mstack_en),
    .wr_en_i_t0(mstack_en_t0)
  );
  paramod85ba01ab5a28334786aba5877c1fe04472f39fbaauxy_ibex_csr  u_mstack_epc_csr (
    .clk_i(clk_i),
    .rd_data_o(mstack_epc_q),
    .rd_data_o_t0(mstack_epc_q_t0),
    .rst_ni(rst_ni),
    .wr_data_i(csr_mepc_o),
    .wr_data_i_t0(csr_mepc_o_t0),
    .wr_en_i(mstack_en),
    .wr_en_i_t0(mstack_en_t0)
  );
  paramod5714e31d82f2b8816750797f158ebea69a089104auxy_ibex_csr  u_mstatus_csr (
    .clk_i(clk_i),
    .rd_data_o(mstatus_q),
    .rd_data_o_t0(mstatus_q_t0),
    .rd_error_o(mstatus_err),
    .rd_error_o_t0(mstatus_err_t0),
    .rst_ni(rst_ni),
    .wr_data_i(mstatus_d),
    .wr_data_i_t0(mstatus_d_t0),
    .wr_en_i(mstatus_en),
    .wr_en_i_t0(mstatus_en_t0)
  );
  paramod85ba01ab5a28334786aba5877c1fe04472f39fbaauxy_ibex_csr  u_mtval_csr (
    .clk_i(clk_i),
    .rd_data_o(mtval_q),
    .rd_data_o_t0(mtval_q_t0),
    .rst_ni(rst_ni),
    .wr_data_i(mtval_d),
    .wr_data_i_t0(mtval_d_t0),
    .wr_en_i(mtval_en),
    .wr_en_i_t0(mtval_en_t0)
  );
  paramod4f46e25470a27719ee9ca03cee1a0827eff766f7auxy_ibex_csr  u_mtvec_csr (
    .clk_i(clk_i),
    .rd_data_o(csr_mtvec_o),
    .rd_data_o_t0(csr_mtvec_o_t0),
    .rd_error_o(mtvec_err),
    .rd_error_o_t0(mtvec_err_t0),
    .rst_ni(rst_ni),
    .wr_data_i(mtvec_d),
    .wr_data_i_t0(mtvec_d_t0),
    .wr_en_i(mtvec_en),
    .wr_en_i_t0(mtvec_en_t0)
  );
  assign { _0000_[31:9], _0000_[5:2] } = { dcsr_d[31:9], dcsr_d[5:2] };
  assign { _0001_[31:9], _0001_[5:2] } = { dcsr_d_t0[31:9], dcsr_d_t0[5:2] };
  assign _0010_[1:0] = mstatus_d[1:0];
  assign _0011_[1:0] = mstatus_d_t0[1:0];
  assign _0022_[8:6] = dcsr_q[8:6];
  assign _0023_[8:6] = dcsr_q_t0[8:6];
  assign csr_mstatus_mie_o = mstatus_q[5];
  assign csr_mstatus_mie_o_t0 = mstatus_q_t0[5];
  assign csr_mstatus_tw_o = mstatus_q[0];
  assign csr_mstatus_tw_o_t0 = mstatus_q_t0[0];
  assign csr_pmp_addr_o = 136'h0000000000000000000000000000000000;
  assign csr_pmp_addr_o_t0 = 136'h0000000000000000000000000000000000;
  assign csr_pmp_cfg_o = 24'h000000;
  assign csr_pmp_cfg_o_t0 = 24'h000000;
  assign csr_pmp_mseccfg_o = 3'h0;
  assign csr_pmp_mseccfg_o_t0 = 3'h0;
  assign data_ind_timing_o = cpuctrl_q[1];
  assign data_ind_timing_o_t0 = cpuctrl_q_t0[1];
  assign debug_ebreakm_o = dcsr_q[15];
  assign debug_ebreakm_o_t0 = dcsr_q_t0[15];
  assign debug_ebreaku_o = dcsr_q[12];
  assign debug_ebreaku_o_t0 = dcsr_q_t0[12];
  assign debug_single_step_o = dcsr_q[2];
  assign debug_single_step_o_t0 = dcsr_q_t0[2];
  assign dummy_instr_en_o = cpuctrl_q[2];
  assign dummy_instr_en_o_t0 = cpuctrl_q_t0[2];
  assign dummy_instr_mask_o = cpuctrl_q[5:3];
  assign dummy_instr_mask_o_t0 = cpuctrl_q_t0[5:3];
  assign dummy_instr_seed_en_o = 1'h0;
  assign dummy_instr_seed_en_o_t0 = 1'h0;
  assign dummy_instr_seed_o = 32'd0;
  assign dummy_instr_seed_o_t0 = 32'd0;
  assign icache_enable_o = cpuctrl_q[0];
  assign icache_enable_o_t0 = cpuctrl_q_t0[0];
  assign { mcountinhibit[31:13], mcountinhibit[1] } = 20'hffffe;
  assign { mcountinhibit_t0[31:13], mcountinhibit_t0[1] } = 20'h00000;
endmodule

module paramodab788080a2d62bee953947d554df7ff9d159e451auxy_ibex_decoder (clk_i, rst_ni, illegal_insn_o, ebrk_insn_o, mret_insn_o, dret_insn_o, ecall_insn_o, wfi_insn_o, jump_set_o, branch_taken_i, icache_inval_o, instr_first_cycle_i, instr_rdata_i, instr_rdata_alu_i, illegal_c_insn_i, imm_a_mux_sel_o, imm_b_mux_sel_o, bt_a_mux_sel_o, bt_b_mux_sel_o, imm_i_type_o, imm_s_type_o
, imm_b_type_o, imm_u_type_o, imm_j_type_o, zimm_rs1_type_o, rf_wdata_sel_o, rf_we_o, rf_raddr_a_o, rf_raddr_b_o, rf_waddr_o, rf_ren_a_o, rf_ren_b_o, alu_operator_o, alu_op_a_mux_sel_o, alu_op_b_mux_sel_o, alu_multicycle_o, mult_en_o, div_en_o, mult_sel_o, div_sel_o, multdiv_operator_o, multdiv_signed_mode_o
, csr_access_o, csr_op_o, data_req_o, data_we_o, data_type_o, data_sign_extension_o, jump_in_dec_o, branch_in_dec_o, instr_rdata_i_t0, alu_multicycle_o_t0, alu_op_a_mux_sel_o_t0, alu_operator_o_t0, branch_in_dec_o_t0, branch_taken_i_t0, bt_b_mux_sel_o_t0, csr_access_o_t0, csr_op_o_t0, data_req_o_t0, data_type_o_t0, div_en_o_t0, div_sel_o_t0
, ebrk_insn_o_t0, ecall_insn_o_t0, icache_inval_o_t0, illegal_insn_o_t0, imm_b_mux_sel_o_t0, imm_i_type_o_t0, imm_j_type_o_t0, imm_s_type_o_t0, imm_u_type_o_t0, instr_rdata_alu_i_t0, jump_set_o_t0, mult_en_o_t0, multdiv_operator_o_t0, multdiv_signed_mode_o_t0, rf_raddr_a_o_t0, rf_ren_a_o_t0, rf_ren_b_o_t0, rf_wdata_sel_o_t0, wfi_insn_o_t0, zimm_rs1_type_o_t0, alu_op_b_mux_sel_o_t0
, rf_we_o_t0, rf_waddr_o_t0, rf_raddr_b_o_t0, mult_sel_o_t0, mret_insn_o_t0, jump_in_dec_o_t0, instr_first_cycle_i_t0, imm_b_type_o_t0, imm_a_mux_sel_o_t0, illegal_c_insn_i_t0, dret_insn_o_t0, data_we_o_t0, data_sign_extension_o_t0, bt_a_mux_sel_o_t0);
  wire [5:0] _0000_;
  wire [5:0] _0001_;
  wire [5:0] _0002_;
  wire [5:0] _0003_;
  wire [5:0] _0004_;
  wire [5:0] _0005_;
  wire _0006_;
  wire _0007_;
  wire [5:0] _0008_;
  wire [5:0] _0009_;
  wire _0010_;
  wire _0011_;
  wire _0012_;
  wire _0013_;
  wire _0014_;
  wire _0015_;
  wire _0016_;
  wire _0017_;
  wire _0018_;
  wire _0019_;
  wire _0020_;
  wire _0021_;
  wire _0022_;
  wire _0023_;
  wire _0024_;
  wire _0025_;
  wire _0026_;
  wire _0027_;
  wire _0028_;
  wire _0029_;
  wire _0030_;
  wire _0031_;
  wire _0032_;
  wire _0033_;
  wire _0034_;
  wire _0035_;
  wire _0036_;
  wire _0037_;
  wire _0038_;
  wire _0039_;
  wire [1:0] _0040_;
  wire [1:0] _0041_;
  wire [1:0] _0042_;
  wire [1:0] _0043_;
  wire _0044_;
  wire _0045_;
  wire _0046_;
  wire _0047_;
  wire _0048_;
  wire _0049_;
  wire _0050_;
  wire _0051_;
  wire _0052_;
  wire _0053_;
  wire _0054_;
  wire _0055_;
  wire _0056_;
  wire _0057_;
  wire _0058_;
  wire _0059_;
  wire _0060_;
  wire _0061_;
  wire _0062_;
  wire _0063_;
  wire [1:0] _0064_;
  wire [1:0] _0065_;
  wire [1:0] _0066_;
  wire [1:0] _0067_;
  wire _0068_;
  wire _0069_;
  wire _0070_;
  wire _0071_;
  wire _0072_;
  wire _0073_;
  wire [1:0] _0074_;
  wire [1:0] _0075_;
  wire _0076_;
  wire _0077_;
  wire _0078_;
  wire _0079_;
  wire _0080_;
  wire _0081_;
  wire _0082_;
  wire _0083_;
  wire _0084_;
  wire _0085_;
  wire _0086_;
  wire _0087_;
  wire _0088_;
  wire _0089_;
  wire [1:0] _0090_;
  wire [1:0] _0091_;
  wire [1:0] _0092_;
  wire [1:0] _0093_;
  wire _0094_;
  wire _0095_;
  wire _0096_;
  wire [1:0] _0097_;
  wire [1:0] _0098_;
  wire _0099_;
  wire [5:0] _0100_;
  wire [5:0] _0101_;
  wire [2:0] _0102_;
  wire [2:0] _0103_;
  wire _0104_;
  wire [2:0] _0105_;
  wire [2:0] _0106_;
  wire [1:0] _0107_;
  wire [1:0] _0108_;
  wire _0109_;
  wire [5:0] _0110_;
  wire [5:0] _0111_;
  wire [2:0] _0112_;
  wire [2:0] _0113_;
  wire _0114_;
  wire _0115_;
  wire [2:0] _0116_;
  wire [2:0] _0117_;
  wire [1:0] _0118_;
  wire [1:0] _0119_;
  wire [5:0] _0120_;
  wire [5:0] _0121_;
  wire _0122_;
  wire _0123_;
  wire [1:0] _0124_;
  wire [1:0] _0125_;
  wire [5:0] _0126_;
  wire [5:0] _0127_;
  wire _0128_;
  wire _0129_;
  wire _0130_;
  wire _0131_;
  wire _0132_;
  wire _0133_;
  wire _0134_;
  wire _0135_;
  wire _0136_;
  wire _0137_;
  wire _0138_;
  wire _0139_;
  wire _0140_;
  wire _0141_;
  wire _0142_;
  wire _0143_;
  wire _0144_;
  wire _0145_;
  wire _0146_;
  wire _0147_;
  wire _0148_;
  wire _0149_;
  wire _0150_;
  wire _0151_;
  wire _0152_;
  wire _0153_;
  wire _0154_;
  wire _0155_;
  wire _0156_;
  wire _0157_;
  wire _0158_;
  wire _0159_;
  wire _0160_;
  wire _0161_;
  wire _0162_;
  wire _0163_;
  wire _0164_;
  wire _0165_;
  wire _0166_;
  wire _0167_;
  wire [1:0] _0168_;
  wire [1:0] _0169_;
  wire [2:0] _0170_;
  wire [1:0] _0171_;
  wire [2:0] _0172_;
  wire [4:0] _0173_;
  wire [5:0] _0174_;
  wire [1:0] _0175_;
  wire [1:0] _0176_;
  wire [2:0] _0177_;
  wire [3:0] _0178_;
  wire [2:0] _0179_;
  wire [3:0] _0180_;
  wire [8:0] _0181_;
  wire [1:0] _0182_;
  wire [1:0] _0183_;
  wire [5:0] _0184_;
  wire [17:0] _0185_;
  wire [5:0] _0186_;
  wire [2:0] _0187_;
  wire [2:0] _0188_;
  wire [1:0] _0189_;
  wire _0190_;
  wire _0191_;
  wire _0192_;
  wire _0193_;
  wire _0194_;
  wire _0195_;
  wire _0196_;
  wire _0197_;
  wire _0198_;
  wire _0199_;
  wire _0200_;
  wire _0201_;
  wire _0202_;
  wire _0203_;
  wire _0204_;
  wire _0205_;
  wire _0206_;
  wire _0207_;
  wire _0208_;
  wire _0209_;
  wire _0210_;
  wire [3:0] _0211_;
  wire [2:0] _0212_;
  wire [2:0] _0213_;
  wire [5:0] _0214_;
  wire [2:0] _0215_;
  wire [5:0] _0216_;
  wire [5:0] _0217_;
  wire [5:0] _0218_;
  wire [5:0] _0219_;
  wire [5:0] _0220_;
  wire [5:0] _0221_;
  wire [5:0] _0222_;
  wire [5:0] _0223_;
  wire [5:0] _0224_;
  wire [5:0] _0225_;
  wire [5:0] _0226_;
  wire [5:0] _0227_;
  wire [5:0] _0228_;
  wire [5:0] _0229_;
  wire [5:0] _0230_;
  wire [5:0] _0231_;
  wire [5:0] _0232_;
  wire [5:0] _0233_;
  wire [5:0] _0234_;
  wire [5:0] _0235_;
  wire [5:0] _0236_;
  wire _0237_;
  wire [1:0] _0238_;
  wire [1:0] _0239_;
  wire [1:0] _0240_;
  wire [1:0] _0241_;
  wire [1:0] _0242_;
  wire [5:0] _0243_;
  wire [5:0] _0244_;
  wire [5:0] _0245_;
  wire [5:0] _0246_;
  wire [5:0] _0247_;
  wire [2:0] _0248_;
  wire [2:0] _0249_;
  wire [2:0] _0250_;
  wire [2:0] _0251_;
  wire [2:0] _0252_;
  wire [2:0] _0253_;
  wire [2:0] _0254_;
  wire [1:0] _0255_;
  wire [1:0] _0256_;
  wire [1:0] _0257_;
  wire [1:0] _0258_;
  wire [1:0] _0259_;
  wire [1:0] _0260_;
  wire [1:0] _0261_;
  wire [1:0] _0262_;
  wire _0263_;
  wire [1:0] _0264_;
  wire _0265_;
  wire _0266_;
  wire _0267_;
  wire _0268_;
  wire _0269_;
  wire [1:0] _0270_;
  wire [4:0] _0271_;
  wire [2:0] _0272_;
  wire [4:0] _0273_;
  wire _0274_;
  wire _0275_;
  wire _0276_;
  wire _0277_;
  wire [2:0] _0278_;
  wire [4:0] _0279_;
  wire [1:0] _0280_;
  wire [1:0] _0281_;
  wire [2:0] _0282_;
  wire [9:0] _0283_;
  wire _0284_;
  wire [5:0] _0285_;
  wire [5:0] _0286_;
  wire [5:0] _0287_;
  wire [2:0] _0288_;
  wire [2:0] _0289_;
  wire [1:0] _0290_;
  wire [5:0] _0291_;
  wire [2:0] _0292_;
  wire [6:0] _0293_;
  wire [1:0] _0294_;
  wire _0295_;
  wire _0296_;
  wire [1:0] _0297_;
  wire _0298_;
  wire _0299_;
  wire [11:0] _0300_;
  wire _0301_;
  wire [1:0] _0302_;
  wire [9:0] _0303_;
  wire _0304_;
  wire [1:0] _0305_;
  wire [1:0] _0306_;
  wire [4:0] _0307_;
  wire _0308_;
  wire [1:0] _0309_;
  wire [5:0] _0310_;
  wire [6:0] _0311_;
  wire [1:0] _0312_;
  wire [1:0] _0313_;
  wire [1:0] _0314_;
  wire [1:0] _0315_;
  wire [2:0] _0316_;
  wire _0317_;
  wire _0318_;
  wire _0319_;
  wire _0320_;
  wire _0321_;
  wire _0322_;
  wire _0323_;
  wire _0324_;
  wire _0325_;
  wire _0326_;
  wire _0327_;
  wire _0328_;
  wire _0329_;
  wire _0330_;
  wire _0331_;
  wire _0332_;
  wire _0333_;
  wire _0334_;
  wire _0335_;
  wire _0336_;
  wire _0337_;
  wire _0338_;
  wire _0339_;
  wire _0340_;
  wire _0341_;
  wire _0342_;
  wire _0343_;
  wire _0344_;
  wire _0345_;
  wire _0346_;
  wire _0347_;
  wire _0348_;
  wire _0349_;
  wire _0350_;
  wire _0351_;
  wire _0352_;
  wire _0353_;
  wire _0354_;
  wire _0355_;
  wire _0356_;
  wire _0357_;
  wire _0358_;
  wire _0359_;
  wire _0360_;
  wire _0361_;
  wire _0362_;
  wire _0363_;
  wire _0364_;
  wire _0365_;
  wire _0366_;
  wire _0367_;
  wire _0368_;
  wire _0369_;
  wire _0370_;
  wire _0371_;
  wire _0372_;
  wire _0373_;
  wire _0374_;
  wire _0375_;
  wire _0376_;
  wire _0377_;
  wire _0378_;
  wire _0379_;
  wire _0380_;
  wire _0381_;
  wire _0382_;
  wire _0383_;
  wire _0384_;
  wire _0385_;
  wire _0386_;
  wire _0387_;
  wire _0388_;
  wire _0389_;
  wire _0390_;
  wire _0391_;
  wire _0392_;
  wire _0393_;
  wire _0394_;
  wire _0395_;
  wire _0396_;
  wire _0397_;
  wire _0398_;
  wire _0399_;
  wire _0400_;
  wire _0401_;
  wire _0402_;
  wire _0403_;
  wire _0404_;
  wire _0405_;
  wire _0406_;
  wire _0407_;
  wire _0408_;
  wire _0409_;
  wire _0410_;
  wire _0411_;
  wire _0412_;
  wire _0413_;
  wire _0414_;
  wire _0415_;
  wire _0416_;
  wire _0417_;
  wire _0418_;
  wire _0419_;
  wire _0420_;
  wire [1:0] _0421_;
  wire [1:0] _0422_;
  wire [2:0] _0423_;
  wire [1:0] _0424_;
  wire [2:0] _0425_;
  wire [4:0] _0426_;
  wire [5:0] _0427_;
  wire [1:0] _0428_;
  wire [1:0] _0429_;
  wire [2:0] _0430_;
  wire [3:0] _0431_;
  wire [2:0] _0432_;
  wire [3:0] _0433_;
  wire [8:0] _0434_;
  wire [1:0] _0435_;
  wire [1:0] _0436_;
  wire [5:0] _0437_;
  wire [17:0] _0438_;
  wire [5:0] _0439_;
  wire [2:0] _0440_;
  wire [2:0] _0441_;
  wire [1:0] _0442_;
  wire _0443_;
  wire _0444_;
  wire _0445_;
  wire _0446_;
  wire _0447_;
  wire _0448_;
  wire _0449_;
  wire _0450_;
  wire _0451_;
  wire _0452_;
  wire _0453_;
  wire _0454_;
  wire _0455_;
  wire _0456_;
  wire _0457_;
  wire _0458_;
  wire _0459_;
  wire _0460_;
  wire _0461_;
  wire _0462_;
  wire _0463_;
  wire _0464_;
  wire _0465_;
  wire _0466_;
  wire _0467_;
  wire _0468_;
  wire _0469_;
  wire _0470_;
  wire _0471_;
  wire _0472_;
  wire _0473_;
  wire _0474_;
  wire _0475_;
  wire _0476_;
  wire _0477_;
  wire _0478_;
  wire [3:0] _0479_;
  wire [2:0] _0480_;
  wire [2:0] _0481_;
  wire [5:0] _0482_;
  wire [2:0] _0483_;
  wire [5:0] _0484_;
  wire [5:0] _0485_;
  wire [5:0] _0486_;
  wire [5:0] _0487_;
  wire [5:0] _0488_;
  wire [5:0] _0489_;
  wire [5:0] _0490_;
  wire [5:0] _0491_;
  wire [5:0] _0492_;
  wire [5:0] _0493_;
  wire [5:0] _0494_;
  wire [5:0] _0495_;
  wire [5:0] _0496_;
  wire [5:0] _0497_;
  wire [5:0] _0498_;
  wire [5:0] _0499_;
  wire [5:0] _0500_;
  wire [5:0] _0501_;
  wire [5:0] _0502_;
  wire [5:0] _0503_;
  wire [5:0] _0504_;
  wire [5:0] _0505_;
  wire [5:0] _0506_;
  wire [5:0] _0507_;
  wire [5:0] _0508_;
  wire [5:0] _0509_;
  wire [5:0] _0510_;
  wire [5:0] _0511_;
  wire [5:0] _0512_;
  wire [5:0] _0513_;
  wire [5:0] _0514_;
  wire [5:0] _0515_;
  wire [5:0] _0516_;
  wire [5:0] _0517_;
  wire [5:0] _0518_;
  wire [5:0] _0519_;
  wire [5:0] _0520_;
  wire [5:0] _0521_;
  wire [5:0] _0522_;
  wire [5:0] _0523_;
  wire [5:0] _0524_;
  wire [5:0] _0525_;
  wire [5:0] _0526_;
  wire [5:0] _0527_;
  wire [5:0] _0528_;
  wire [5:0] _0529_;
  wire [5:0] _0530_;
  wire [5:0] _0531_;
  wire [5:0] _0532_;
  wire [5:0] _0533_;
  wire [5:0] _0534_;
  wire [5:0] _0535_;
  wire [5:0] _0536_;
  wire [5:0] _0537_;
  wire [5:0] _0538_;
  wire [5:0] _0539_;
  wire [5:0] _0540_;
  wire [5:0] _0541_;
  wire [5:0] _0542_;
  wire [5:0] _0543_;
  wire [5:0] _0544_;
  wire [5:0] _0545_;
  wire [5:0] _0546_;
  wire [5:0] _0547_;
  wire _0548_;
  wire _0549_;
  wire _0550_;
  wire _0551_;
  wire _0552_;
  wire _0553_;
  wire _0554_;
  wire [1:0] _0555_;
  wire [1:0] _0556_;
  wire [1:0] _0557_;
  wire [1:0] _0558_;
  wire [1:0] _0559_;
  wire [1:0] _0560_;
  wire [1:0] _0561_;
  wire [1:0] _0562_;
  wire [1:0] _0563_;
  wire [1:0] _0564_;
  wire [1:0] _0565_;
  wire [1:0] _0566_;
  wire [1:0] _0567_;
  wire [1:0] _0568_;
  wire [1:0] _0569_;
  wire [5:0] _0570_;
  wire [5:0] _0571_;
  wire [5:0] _0572_;
  wire [5:0] _0573_;
  wire [5:0] _0574_;
  wire [5:0] _0575_;
  wire [5:0] _0576_;
  wire [5:0] _0577_;
  wire [5:0] _0578_;
  wire [5:0] _0579_;
  wire [5:0] _0580_;
  wire [5:0] _0581_;
  wire [5:0] _0582_;
  wire [5:0] _0583_;
  wire [5:0] _0584_;
  wire [2:0] _0585_;
  wire [2:0] _0586_;
  wire [2:0] _0587_;
  wire [2:0] _0588_;
  wire [2:0] _0589_;
  wire [2:0] _0590_;
  wire [2:0] _0591_;
  wire [2:0] _0592_;
  wire [2:0] _0593_;
  wire [2:0] _0594_;
  wire [2:0] _0595_;
  wire [2:0] _0596_;
  wire [2:0] _0597_;
  wire [2:0] _0598_;
  wire [2:0] _0599_;
  wire [2:0] _0600_;
  wire [2:0] _0601_;
  wire [2:0] _0602_;
  wire [2:0] _0603_;
  wire [2:0] _0604_;
  wire [2:0] _0605_;
  wire [1:0] _0606_;
  wire [1:0] _0607_;
  wire [1:0] _0608_;
  wire [1:0] _0609_;
  wire [1:0] _0610_;
  wire [1:0] _0611_;
  wire [1:0] _0612_;
  wire [1:0] _0613_;
  wire [1:0] _0614_;
  wire [1:0] _0615_;
  wire [1:0] _0616_;
  wire [1:0] _0617_;
  wire [1:0] _0618_;
  wire [1:0] _0619_;
  wire [1:0] _0620_;
  wire [1:0] _0621_;
  wire [1:0] _0622_;
  wire [1:0] _0623_;
  wire [1:0] _0624_;
  wire [1:0] _0625_;
  wire [1:0] _0626_;
  wire [1:0] _0627_;
  wire [1:0] _0628_;
  wire [1:0] _0629_;
  wire _0630_;
  wire _0631_;
  wire _0632_;
  wire _0633_;
  wire _0634_;
  wire _0635_;
  wire _0636_;
  wire _0637_;
  wire [1:0] _0638_;
  wire [1:0] _0639_;
  wire [1:0] _0640_;
  wire [1:0] _0641_;
  wire [1:0] _0642_;
  wire _0643_;
  wire _0644_;
  wire _0645_;
  wire _0646_;
  wire _0647_;
  wire _0648_;
  wire _0649_;
  wire _0650_;
  wire _0651_;
  wire _0652_;
  wire _0653_;
  wire _0654_;
  wire _0655_;
  wire _0656_;
  wire _0657_;
  wire _0658_;
  wire _0659_;
  wire _0660_;
  wire _0661_;
  wire _0662_;
  wire _0663_;
  wire _0664_;
  wire _0665_;
  wire _0666_;
  wire _0667_;
  wire _0668_;
  wire _0669_;
  wire _0670_;
  wire _0671_;
  wire _0672_;
  wire _0673_;
  wire _0674_;
  wire _0675_;
  wire _0676_;
  wire _0677_;
  wire _0678_;
  wire _0679_;
  wire _0680_;
  wire _0681_;
  wire [1:0] _0682_;
  wire [1:0] _0683_;
  wire [1:0] _0684_;
  wire [4:0] _0685_;
  wire [2:0] _0686_;
  wire [2:0] _0687_;
  wire [4:0] _0688_;
  wire [4:0] _0689_;
  wire _0690_;
  wire _0691_;
  wire _0692_;
  wire _0693_;
  wire _0694_;
  wire _0695_;
  wire _0696_;
  wire _0697_;
  wire _0698_;
  wire [2:0] _0699_;
  wire [4:0] _0700_;
  wire [1:0] _0701_;
  wire [1:0] _0702_;
  wire [1:0] _0703_;
  wire [1:0] _0704_;
  wire [1:0] _0705_;
  wire [1:0] _0706_;
  wire [1:0] _0707_;
  wire [1:0] _0708_;
  wire [5:0] _0709_;
  wire [2:0] _0710_;
  wire [2:0] _0711_;
  wire [2:0] _0712_;
  wire [9:0] _0713_;
  wire [9:0] _0714_;
  wire [9:0] _0715_;
  wire [9:0] _0716_;
  wire [9:0] _0717_;
  wire [9:0] _0718_;
  wire [9:0] _0719_;
  wire [9:0] _0720_;
  wire [9:0] _0721_;
  wire [9:0] _0722_;
  wire [9:0] _0723_;
  wire [9:0] _0724_;
  wire [9:0] _0725_;
  wire [9:0] _0726_;
  wire [9:0] _0727_;
  wire [9:0] _0728_;
  wire [9:0] _0729_;
  wire _0730_;
  wire _0731_;
  wire _0732_;
  wire _0733_;
  wire [5:0] _0734_;
  wire [5:0] _0735_;
  wire [5:0] _0736_;
  wire [5:0] _0737_;
  wire [5:0] _0738_;
  wire [5:0] _0739_;
  wire [5:0] _0740_;
  wire [5:0] _0741_;
  wire [5:0] _0742_;
  wire [2:0] _0743_;
  wire [2:0] _0744_;
  wire [2:0] _0745_;
  wire [2:0] _0746_;
  wire [2:0] _0747_;
  wire [2:0] _0748_;
  wire [1:0] _0749_;
  wire [1:0] _0750_;
  wire [1:0] _0751_;
  wire [5:0] _0752_;
  wire [5:0] _0753_;
  wire [5:0] _0754_;
  wire [2:0] _0755_;
  wire [2:0] _0756_;
  wire [2:0] _0757_;
  wire [2:0] _0758_;
  wire [2:0] _0759_;
  wire [2:0] _0760_;
  wire [2:0] _0761_;
  wire [2:0] _0762_;
  wire [6:0] _0763_;
  wire [6:0] _0764_;
  wire [6:0] _0765_;
  wire [6:0] _0766_;
  wire [6:0] _0767_;
  wire [6:0] _0768_;
  wire [1:0] _0769_;
  wire [1:0] _0770_;
  wire [1:0] _0771_;
  wire [6:0] _0772_;
  wire [6:0] _0773_;
  wire [6:0] _0774_;
  wire [6:0] _0775_;
  wire _0776_;
  wire _0777_;
  wire _0778_;
  wire _0779_;
  wire [6:0] _0780_;
  wire _0781_;
  wire _0782_;
  wire [6:0] _0783_;
  wire _0784_;
  wire _0785_;
  wire _0786_;
  wire _0787_;
  wire _0788_;
  wire _0789_;
  wire _0790_;
  wire _0791_;
  wire _0792_;
  wire _0793_;
  wire _0794_;
  wire _0795_;
  wire _0796_;
  wire _0797_;
  wire _0798_;
  wire _0799_;
  wire [1:0] _0800_;
  wire [1:0] _0801_;
  wire _0802_;
  wire _0803_;
  wire [11:0] _0804_;
  wire [11:0] _0805_;
  wire [11:0] _0806_;
  wire [11:0] _0807_;
  wire [11:0] _0808_;
  wire _0809_;
  wire _0810_;
  wire _0811_;
  wire _0812_;
  wire _0813_;
  wire _0814_;
  wire _0815_;
  wire _0816_;
  wire _0817_;
  wire _0818_;
  wire _0819_;
  wire _0820_;
  wire _0821_;
  wire _0822_;
  wire _0823_;
  wire [1:0] _0824_;
  wire [1:0] _0825_;
  wire [1:0] _0826_;
  wire _0827_;
  wire _0828_;
  wire [9:0] _0829_;
  wire [9:0] _0830_;
  wire [9:0] _0831_;
  wire [9:0] _0832_;
  wire [9:0] _0833_;
  wire [9:0] _0834_;
  wire [9:0] _0835_;
  wire [9:0] _0836_;
  wire [9:0] _0837_;
  wire [9:0] _0838_;
  wire [9:0] _0839_;
  wire [9:0] _0840_;
  wire [9:0] _0841_;
  wire [9:0] _0842_;
  wire [9:0] _0843_;
  wire [9:0] _0844_;
  wire [9:0] _0845_;
  wire [9:0] _0846_;
  wire _0847_;
  wire _0848_;
  wire [1:0] _0849_;
  wire [1:0] _0850_;
  wire [1:0] _0851_;
  wire [1:0] _0852_;
  wire [1:0] _0853_;
  wire _0854_;
  wire _0855_;
  wire [1:0] _0856_;
  wire [4:0] _0857_;
  wire [4:0] _0858_;
  wire _0859_;
  wire _0860_;
  wire [1:0] _0861_;
  wire _0862_;
  wire _0863_;
  wire _0864_;
  wire _0865_;
  wire [1:0] _0866_;
  wire [1:0] _0867_;
  wire [5:0] _0868_;
  wire [2:0] _0869_;
  wire [2:0] _0870_;
  wire [2:0] _0871_;
  wire [2:0] _0872_;
  wire [2:0] _0873_;
  wire [6:0] _0874_;
  wire [6:0] _0875_;
  wire [6:0] _0876_;
  wire [6:0] _0877_;
  wire [6:0] _0878_;
  wire _0879_;
  wire _0880_;
  wire [1:0] _0881_;
  wire [1:0] _0882_;
  wire [1:0] _0883_;
  wire [1:0] _0884_;
  wire [1:0] _0885_;
  wire [1:0] _0886_;
  wire [1:0] _0887_;
  wire [1:0] _0888_;
  wire _0889_;
  wire _0890_;
  wire _0891_;
  wire _0892_;
  wire _0893_;
  wire _0894_;
  wire _0895_;
  wire _0896_;
  wire _0897_;
  wire _0898_;
  wire _0899_;
  wire [6:0] _0900_;
  wire [6:0] _0901_;
  wire [6:0] _0902_;
  wire [6:0] _0903_;
  wire [6:0] _0904_;
  wire [6:0] _0905_;
  wire [6:0] _0906_;
  wire _0907_;
  wire [1:0] _0908_;
  wire [1:0] _0909_;
  wire [1:0] _0910_;
  wire [1:0] _0911_;
  wire [1:0] _0912_;
  wire [1:0] _0913_;
  wire _0914_;
  wire [2:0] _0915_;
  wire [2:0] _0916_;
  wire [2:0] _0917_;
  wire _0918_;
  wire _0919_;
  wire _0920_;
  wire _0921_;
  wire _0922_;
  wire _0923_;
  wire _0924_;
  wire _0925_;
  wire _0926_;
  wire _0927_;
  wire _0928_;
  wire _0929_;
  wire _0930_;
  wire _0931_;
  wire _0932_;
  wire _0933_;
  wire _0934_;
  wire _0935_;
  wire _0936_;
  wire _0937_;
  wire _0938_;
  wire _0939_;
  wire _0940_;
  wire _0941_;
  wire _0942_;
  wire _0943_;
  wire _0944_;
  wire _0945_;
  wire _0946_;
  wire _0947_;
  wire _0948_;
  wire _0949_;
  wire _0950_;
  wire _0951_;
  wire _0952_;
  wire _0953_;
  wire _0954_;
  wire _0955_;
  wire _0956_;
  wire _0957_;
  wire [5:0] _0958_;
  wire [5:0] _0959_;
  wire [5:0] _0960_;
  wire [5:0] _0961_;
  wire [5:0] _0962_;
  wire [5:0] _0963_;
  wire [5:0] _0964_;
  wire [5:0] _0965_;
  wire [5:0] _0966_;
  wire [5:0] _0967_;
  wire [5:0] _0968_;
  wire [5:0] _0969_;
  wire [5:0] _0970_;
  wire [5:0] _0971_;
  wire [5:0] _0972_;
  wire [5:0] _0973_;
  wire [5:0] _0974_;
  wire [5:0] _0975_;
  wire [5:0] _0976_;
  wire [5:0] _0977_;
  wire [5:0] _0978_;
  wire [5:0] _0979_;
  wire [5:0] _0980_;
  wire [5:0] _0981_;
  wire [5:0] _0982_;
  wire [5:0] _0983_;
  wire [5:0] _0984_;
  wire [5:0] _0985_;
  wire [5:0] _0986_;
  wire [5:0] _0987_;
  wire [5:0] _0988_;
  wire [5:0] _0989_;
  wire [5:0] _0990_;
  wire [5:0] _0991_;
  wire [5:0] _0992_;
  wire [5:0] _0993_;
  wire [5:0] _0994_;
  wire [5:0] _0995_;
  wire [5:0] _0996_;
  wire [5:0] _0997_;
  wire [5:0] _0998_;
  wire [5:0] _0999_;
  wire [5:0] _1000_;
  wire [5:0] _1001_;
  wire [5:0] _1002_;
  wire [5:0] _1003_;
  wire [5:0] _1004_;
  wire [5:0] _1005_;
  wire [5:0] _1006_;
  wire [5:0] _1007_;
  wire [5:0] _1008_;
  wire [5:0] _1009_;
  wire [5:0] _1010_;
  wire [5:0] _1011_;
  wire [5:0] _1012_;
  wire [5:0] _1013_;
  wire [5:0] _1014_;
  wire [5:0] _1015_;
  wire [5:0] _1016_;
  wire [5:0] _1017_;
  wire [5:0] _1018_;
  wire _1019_;
  wire _1020_;
  wire _1021_;
  wire _1022_;
  wire _1023_;
  wire _1024_;
  wire [1:0] _1025_;
  wire [1:0] _1026_;
  wire [1:0] _1027_;
  wire [1:0] _1028_;
  wire [1:0] _1029_;
  wire [1:0] _1030_;
  wire [1:0] _1031_;
  wire [1:0] _1032_;
  wire [1:0] _1033_;
  wire [1:0] _1034_;
  wire [1:0] _1035_;
  wire [1:0] _1036_;
  wire [1:0] _1037_;
  wire [1:0] _1038_;
  wire [1:0] _1039_;
  wire [5:0] _1040_;
  wire [5:0] _1041_;
  wire [5:0] _1042_;
  wire [5:0] _1043_;
  wire [5:0] _1044_;
  wire [5:0] _1045_;
  wire [5:0] _1046_;
  wire [5:0] _1047_;
  wire [5:0] _1048_;
  wire [5:0] _1049_;
  wire [5:0] _1050_;
  wire [5:0] _1051_;
  wire [5:0] _1052_;
  wire [5:0] _1053_;
  wire [5:0] _1054_;
  wire [2:0] _1055_;
  wire [2:0] _1056_;
  wire [2:0] _1057_;
  wire [2:0] _1058_;
  wire [2:0] _1059_;
  wire [2:0] _1060_;
  wire [2:0] _1061_;
  wire [2:0] _1062_;
  wire [2:0] _1063_;
  wire [2:0] _1064_;
  wire [2:0] _1065_;
  wire [2:0] _1066_;
  wire [2:0] _1067_;
  wire [2:0] _1068_;
  wire [2:0] _1069_;
  wire [2:0] _1070_;
  wire [2:0] _1071_;
  wire [2:0] _1072_;
  wire [2:0] _1073_;
  wire [2:0] _1074_;
  wire [2:0] _1075_;
  wire [1:0] _1076_;
  wire [1:0] _1077_;
  wire [1:0] _1078_;
  wire [1:0] _1079_;
  wire [1:0] _1080_;
  wire [1:0] _1081_;
  wire [1:0] _1082_;
  wire [1:0] _1083_;
  wire [1:0] _1084_;
  wire [1:0] _1085_;
  wire [1:0] _1086_;
  wire [1:0] _1087_;
  wire [1:0] _1088_;
  wire [1:0] _1089_;
  wire [1:0] _1090_;
  wire [1:0] _1091_;
  wire [1:0] _1092_;
  wire [1:0] _1093_;
  wire [1:0] _1094_;
  wire [1:0] _1095_;
  wire [1:0] _1096_;
  wire [1:0] _1097_;
  wire [1:0] _1098_;
  wire [1:0] _1099_;
  wire _1100_;
  wire _1101_;
  wire _1102_;
  wire _1103_;
  wire _1104_;
  wire _1105_;
  wire _1106_;
  wire [1:0] _1107_;
  wire [1:0] _1108_;
  wire [1:0] _1109_;
  wire [1:0] _1110_;
  wire _1111_;
  wire _1112_;
  wire _1113_;
  wire _1114_;
  wire _1115_;
  wire _1116_;
  wire _1117_;
  wire _1118_;
  wire _1119_;
  wire _1120_;
  wire _1121_;
  wire _1122_;
  wire _1123_;
  wire _1124_;
  wire _1125_;
  wire _1126_;
  wire _1127_;
  wire _1128_;
  wire _1129_;
  wire _1130_;
  wire _1131_;
  wire _1132_;
  wire _1133_;
  wire _1134_;
  wire _1135_;
  wire _1136_;
  wire _1137_;
  wire _1138_;
  wire _1139_;
  wire _1140_;
  wire _1141_;
  wire _1142_;
  wire _1143_;
  wire [1:0] _1144_;
  wire [1:0] _1145_;
  wire [1:0] _1146_;
  wire [1:0] _1147_;
  wire [1:0] _1148_;
  wire [1:0] _1149_;
  wire [1:0] _1150_;
  wire [2:0] _1151_;
  wire [2:0] _1152_;
  wire [2:0] _1153_;
  wire _1154_;
  wire [5:0] _1155_;
  wire [5:0] _1156_;
  wire [5:0] _1157_;
  wire [5:0] _1158_;
  wire [5:0] _1159_;
  wire [5:0] _1160_;
  wire [5:0] _1161_;
  wire [5:0] _1162_;
  wire [5:0] _1163_;
  wire [2:0] _1164_;
  wire [2:0] _1165_;
  wire [2:0] _1166_;
  wire [1:0] _1167_;
  wire [1:0] _1168_;
  wire [1:0] _1169_;
  wire [5:0] _1170_;
  wire [5:0] _1171_;
  wire [5:0] _1172_;
  wire [2:0] _1173_;
  wire [2:0] _1174_;
  wire [2:0] _1175_;
  wire [1:0] _1176_;
  wire [1:0] _1177_;
  wire [1:0] _1178_;
  wire _1179_;
  wire _1180_;
  wire _1181_;
  wire _1182_;
  wire _1183_;
  wire _1184_;
  wire _1185_;
  wire [1:0] _1186_;
  wire [1:0] _1187_;
  wire [1:0] _1188_;
  wire _1189_;
  wire [1:0] _1190_;
  wire [1:0] _1191_;
  wire [1:0] _1192_;
  wire [1:0] _1193_;
  wire _1194_;
  wire _1195_;
  wire _1196_;
  wire _1197_;
  wire [1:0] _1198_;
  wire [1:0] _1199_;
  wire [1:0] _1200_;
  wire [1:0] _1201_;
  wire [1:0] _1202_;
  wire [1:0] _1203_;
  wire [1:0] _1204_;
  wire [1:0] _1205_;
  wire [1:0] _1206_;
  wire [1:0] _1207_;
  wire [1:0] _1208_;
  wire [1:0] _1209_;
  wire [1:0] _1210_;
  wire [2:0] _1211_;
  wire [2:0] _1212_;
  wire [2:0] _1213_;
  wire [5:0] _1214_;
  wire [5:0] _1215_;
  wire [5:0] _1216_;
  wire [5:0] _1217_;
  wire [5:0] _1218_;
  wire [5:0] _1219_;
  wire [5:0] _1220_;
  wire [5:0] _1221_;
  wire [5:0] _1222_;
  wire [5:0] _1223_;
  wire [5:0] _1224_;
  wire [5:0] _1225_;
  wire _1226_;
  wire [1:0] _1227_;
  wire [1:0] _1228_;
  wire [1:0] _1229_;
  wire [1:0] _1230_;
  wire [5:0] _1231_;
  wire [5:0] _1232_;
  wire [5:0] _1233_;
  wire [5:0] _1234_;
  wire [5:0] _1235_;
  wire [2:0] _1236_;
  wire [2:0] _1237_;
  wire [2:0] _1238_;
  wire [2:0] _1239_;
  wire [2:0] _1240_;
  wire [1:0] _1241_;
  wire [1:0] _1242_;
  wire [1:0] _1243_;
  wire _1244_;
  wire _1245_;
  wire [1:0] _1246_;
  wire _1247_;
  wire _1248_;
  wire _1249_;
  wire _1250_;
  wire _1251_;
  wire _1252_;
  wire _1253_;
  wire _1254_;
  wire _1255_;
  wire _1256_;
  wire _1257_;
  wire [5:0] _1258_;
  wire [5:0] _1259_;
  wire _1260_;
  wire _1261_;
  wire _1262_;
  wire _1263_;
  wire _1264_;
  wire _1265_;
  wire _1266_;
  wire _1267_;
  wire _1268_;
  wire _1269_;
  wire _1270_;
  wire _1271_;
  wire _1272_;
  wire _1273_;
  wire _1274_;
  wire _1275_;
  wire _1276_;
  wire _1277_;
  wire _1278_;
  wire _1279_;
  wire _1280_;
  wire _1281_;
  wire _1282_;
  wire _1283_;
  wire _1284_;
  wire _1285_;
  wire _1286_;
  wire _1287_;
  wire _1288_;
  wire _1289_;
  wire _1290_;
  wire _1291_;
  wire _1292_;
  wire _1293_;
  wire _1294_;
  wire _1295_;
  wire _1296_;
  wire _1297_;
  wire _1298_;
  wire _1299_;
  wire _1300_;
  wire _1301_;
  wire _1302_;
  wire _1303_;
  wire _1304_;
  wire _1305_;
  wire _1306_;
  wire _1307_;
  wire _1308_;
  wire _1309_;
  wire _1310_;
  wire _1311_;
  wire _1312_;
  wire _1313_;
  wire _1314_;
  wire _1315_;
  wire _1316_;
  wire _1317_;
  wire _1318_;
  wire _1319_;
  wire _1320_;
  wire _1321_;
  wire _1322_;
  wire _1323_;
  wire _1324_;
  wire _1325_;
  wire _1326_;
  wire _1327_;
  wire _1328_;
  wire _1329_;
  wire _1330_;
  wire _1331_;
  wire _1332_;
  wire _1333_;
  wire _1334_;
  wire _1335_;
  wire _1336_;
  wire _1337_;
  wire _1338_;
  wire _1339_;
  wire [5:0] _1340_;
  wire [5:0] _1341_;
  wire [5:0] _1342_;
  wire [5:0] _1343_;
  wire [5:0] _1344_;
  wire [5:0] _1345_;
  wire [5:0] _1346_;
  wire [5:0] _1347_;
  wire [5:0] _1348_;
  wire [5:0] _1349_;
  wire [5:0] _1350_;
  wire [5:0] _1351_;
  wire [5:0] _1352_;
  wire [5:0] _1353_;
  wire [5:0] _1354_;
  wire [5:0] _1355_;
  wire [5:0] _1356_;
  wire [5:0] _1357_;
  wire [5:0] _1358_;
  wire [5:0] _1359_;
  wire [5:0] _1360_;
  wire [5:0] _1361_;
  wire [5:0] _1362_;
  wire [5:0] _1363_;
  wire [5:0] _1364_;
  wire [5:0] _1365_;
  wire [5:0] _1366_;
  wire [5:0] _1367_;
  wire [5:0] _1368_;
  wire [5:0] _1369_;
  wire [5:0] _1370_;
  wire [5:0] _1371_;
  wire [5:0] _1372_;
  wire [5:0] _1373_;
  wire [5:0] _1374_;
  wire [5:0] _1375_;
  wire [5:0] _1376_;
  wire [5:0] _1377_;
  wire _1378_;
  wire _1379_;
  wire _1380_;
  wire _1381_;
  wire [1:0] _1382_;
  wire [1:0] _1383_;
  wire [1:0] _1384_;
  wire [1:0] _1385_;
  wire [1:0] _1386_;
  wire [1:0] _1387_;
  wire [1:0] _1388_;
  wire [1:0] _1389_;
  wire [5:0] _1390_;
  wire [5:0] _1391_;
  wire [5:0] _1392_;
  wire [5:0] _1393_;
  wire [5:0] _1394_;
  wire [5:0] _1395_;
  wire [5:0] _1396_;
  wire [2:0] _1397_;
  wire [2:0] _1398_;
  wire [2:0] _1399_;
  wire [2:0] _1400_;
  wire [2:0] _1401_;
  wire [2:0] _1402_;
  wire [2:0] _1403_;
  wire [2:0] _1404_;
  wire [2:0] _1405_;
  wire [2:0] _1406_;
  wire [1:0] _1407_;
  wire [1:0] _1408_;
  wire [1:0] _1409_;
  wire [1:0] _1410_;
  wire [1:0] _1411_;
  wire [1:0] _1412_;
  wire [1:0] _1413_;
  wire [1:0] _1414_;
  wire [1:0] _1415_;
  wire [1:0] _1416_;
  wire _1417_;
  wire _1418_;
  wire _1419_;
  wire [1:0] _1420_;
  wire [1:0] _1421_;
  wire _1422_;
  wire _1423_;
  wire _1424_;
  wire _1425_;
  wire _1426_;
  wire _1427_;
  wire _1428_;
  wire _1429_;
  wire _1430_;
  wire _1431_;
  wire _1432_;
  wire _1433_;
  wire _1434_;
  wire _1435_;
  wire _1436_;
  wire _1437_;
  wire _1438_;
  wire _1439_;
  wire _1440_;
  wire _1441_;
  wire _1442_;
  wire _1443_;
  wire _1444_;
  wire _1445_;
  wire _1446_;
  wire _1447_;
  wire _1448_;
  wire _1449_;
  wire _1450_;
  wire _1451_;
  wire _1452_;
  wire _1453_;
  wire _1454_;
  wire _1455_;
  wire _1456_;
  wire _1457_;
  wire _1458_;
  wire _1459_;
  wire _1460_;
  wire _1461_;
  wire _1462_;
  wire _1463_;
  wire _1464_;
  wire _1465_;
  wire _1466_;
  wire _1467_;
  wire _1468_;
  wire _1469_;
  wire _1470_;
  wire _1471_;
  wire _1472_;
  wire _1473_;
  wire _1474_;
  wire _1475_;
  wire _1476_;
  wire _1477_;
  wire _1478_;
  wire _1479_;
  wire _1480_;
  wire _1481_;
  wire _1482_;
  wire _1483_;
  wire _1484_;
  wire _1485_;
  wire _1486_;
  wire _1487_;
  wire _1488_;
  wire _1489_;
  wire _1490_;
  wire _1491_;
  wire _1492_;
  wire _1493_;
  wire _1494_;
  wire _1495_;
  wire _1496_;
  wire _1497_;
  wire _1498_;
  wire _1499_;
  wire _1500_;
  wire _1501_;
  wire _1502_;
  wire _1503_;
  wire _1504_;
  wire _1505_;
  wire _1506_;
  wire _1507_;
  wire _1508_;
  wire _1509_;
  wire _1510_;
  wire _1511_;
  wire _1512_;
  wire _1513_;
  wire _1514_;
  wire _1515_;
  wire _1516_;
  wire _1517_;
  wire _1518_;
  wire _1519_;
  wire _1520_;
  wire _1521_;
  wire _1522_;
  wire _1523_;
  wire _1524_;
  wire _1525_;
  wire _1526_;
  wire _1527_;
  wire _1528_;
  wire _1529_;
  wire _1530_;
  wire _1531_;
  wire _1532_;
  wire _1533_;
  wire _1534_;
  wire _1535_;
  wire _1536_;
  wire _1537_;
  wire _1538_;
  wire _1539_;
  wire _1540_;
  wire _1541_;
  wire _1542_;
  wire _1543_;
  wire _1544_;
  wire _1545_;
  wire _1546_;
  wire _1547_;
  wire _1548_;
  wire _1549_;
  wire _1550_;
  wire _1551_;
  wire _1552_;
  wire _1553_;
  wire _1554_;
  wire _1555_;
  wire _1556_;
  wire _1557_;
  wire _1558_;
  wire _1559_;
  wire _1560_;
  wire _1561_;
  wire _1562_;
  wire _1563_;
  wire _1564_;
  wire _1565_;
  wire _1566_;
  wire _1567_;
  wire _1568_;
  wire [9:0] _1569_;
  wire [9:0] _1570_;
  wire _1571_;
  wire _1572_;
  wire _1573_;
  wire _1574_;
  wire _1575_;
  wire _1576_;
  wire [1:0] _1577_;
  wire [1:0] _1578_;
  wire _1579_;
  wire _1580_;
  wire [5:0] _1581_;
  wire [5:0] _1582_;
  wire _1583_;
  wire _1584_;
  wire _1585_;
  wire _1586_;
  wire _1587_;
  wire _1588_;
  wire _1589_;
  wire _1590_;
  wire _1591_;
  wire _1592_;
  wire _1593_;
  wire _1594_;
  wire _1595_;
  wire _1596_;
  wire _1597_;
  wire _1598_;
  output alu_multicycle_o;
  wire alu_multicycle_o;
  output alu_multicycle_o_t0;
  wire alu_multicycle_o_t0;
  output [1:0] alu_op_a_mux_sel_o;
  wire [1:0] alu_op_a_mux_sel_o;
  output [1:0] alu_op_a_mux_sel_o_t0;
  wire [1:0] alu_op_a_mux_sel_o_t0;
  output alu_op_b_mux_sel_o;
  wire alu_op_b_mux_sel_o;
  output alu_op_b_mux_sel_o_t0;
  wire alu_op_b_mux_sel_o_t0;
  output [5:0] alu_operator_o;
  wire [5:0] alu_operator_o;
  output [5:0] alu_operator_o_t0;
  wire [5:0] alu_operator_o_t0;
  output branch_in_dec_o;
  wire branch_in_dec_o;
  output branch_in_dec_o_t0;
  wire branch_in_dec_o_t0;
  input branch_taken_i;
  wire branch_taken_i;
  input branch_taken_i_t0;
  wire branch_taken_i_t0;
  output [1:0] bt_a_mux_sel_o;
  wire [1:0] bt_a_mux_sel_o;
  output [1:0] bt_a_mux_sel_o_t0;
  wire [1:0] bt_a_mux_sel_o_t0;
  output [2:0] bt_b_mux_sel_o;
  wire [2:0] bt_b_mux_sel_o;
  output [2:0] bt_b_mux_sel_o_t0;
  wire [2:0] bt_b_mux_sel_o_t0;
  input clk_i;
  wire clk_i;
  output csr_access_o;
  wire csr_access_o;
  output csr_access_o_t0;
  wire csr_access_o_t0;
  wire [1:0] csr_op;
  output [1:0] csr_op_o;
  wire [1:0] csr_op_o;
  output [1:0] csr_op_o_t0;
  wire [1:0] csr_op_o_t0;
  wire [1:0] csr_op_t0;
  output data_req_o;
  wire data_req_o;
  output data_req_o_t0;
  wire data_req_o_t0;
  output data_sign_extension_o;
  wire data_sign_extension_o;
  output data_sign_extension_o_t0;
  wire data_sign_extension_o_t0;
  output [1:0] data_type_o;
  wire [1:0] data_type_o;
  output [1:0] data_type_o_t0;
  wire [1:0] data_type_o_t0;
  output data_we_o;
  wire data_we_o;
  output data_we_o_t0;
  wire data_we_o_t0;
  output div_en_o;
  wire div_en_o;
  output div_en_o_t0;
  wire div_en_o_t0;
  output div_sel_o;
  wire div_sel_o;
  output div_sel_o_t0;
  wire div_sel_o_t0;
  output dret_insn_o;
  wire dret_insn_o;
  output dret_insn_o_t0;
  wire dret_insn_o_t0;
  output ebrk_insn_o;
  wire ebrk_insn_o;
  output ebrk_insn_o_t0;
  wire ebrk_insn_o_t0;
  output ecall_insn_o;
  wire ecall_insn_o;
  output ecall_insn_o_t0;
  wire ecall_insn_o_t0;
  output icache_inval_o;
  wire icache_inval_o;
  output icache_inval_o_t0;
  wire icache_inval_o_t0;
  input illegal_c_insn_i;
  wire illegal_c_insn_i;
  input illegal_c_insn_i_t0;
  wire illegal_c_insn_i_t0;
  output illegal_insn_o;
  wire illegal_insn_o;
  output illegal_insn_o_t0;
  wire illegal_insn_o_t0;
  output imm_a_mux_sel_o;
  wire imm_a_mux_sel_o;
  output imm_a_mux_sel_o_t0;
  wire imm_a_mux_sel_o_t0;
  output [2:0] imm_b_mux_sel_o;
  wire [2:0] imm_b_mux_sel_o;
  output [2:0] imm_b_mux_sel_o_t0;
  wire [2:0] imm_b_mux_sel_o_t0;
  output [31:0] imm_b_type_o;
  wire [31:0] imm_b_type_o;
  output [31:0] imm_b_type_o_t0;
  wire [31:0] imm_b_type_o_t0;
  output [31:0] imm_i_type_o;
  wire [31:0] imm_i_type_o;
  output [31:0] imm_i_type_o_t0;
  wire [31:0] imm_i_type_o_t0;
  output [31:0] imm_j_type_o;
  wire [31:0] imm_j_type_o;
  output [31:0] imm_j_type_o_t0;
  wire [31:0] imm_j_type_o_t0;
  output [31:0] imm_s_type_o;
  wire [31:0] imm_s_type_o;
  output [31:0] imm_s_type_o_t0;
  wire [31:0] imm_s_type_o_t0;
  output [31:0] imm_u_type_o;
  wire [31:0] imm_u_type_o;
  output [31:0] imm_u_type_o_t0;
  wire [31:0] imm_u_type_o_t0;
  input instr_first_cycle_i;
  wire instr_first_cycle_i;
  input instr_first_cycle_i_t0;
  wire instr_first_cycle_i_t0;
  input [31:0] instr_rdata_alu_i;
  wire [31:0] instr_rdata_alu_i;
  input [31:0] instr_rdata_alu_i_t0;
  wire [31:0] instr_rdata_alu_i_t0;
  input [31:0] instr_rdata_i;
  wire [31:0] instr_rdata_i;
  input [31:0] instr_rdata_i_t0;
  wire [31:0] instr_rdata_i_t0;
  output jump_in_dec_o;
  wire jump_in_dec_o;
  output jump_in_dec_o_t0;
  wire jump_in_dec_o_t0;
  output jump_set_o;
  wire jump_set_o;
  output jump_set_o_t0;
  wire jump_set_o_t0;
  output mret_insn_o;
  wire mret_insn_o;
  output mret_insn_o_t0;
  wire mret_insn_o_t0;
  output mult_en_o;
  wire mult_en_o;
  output mult_en_o_t0;
  wire mult_en_o_t0;
  output mult_sel_o;
  wire mult_sel_o;
  output mult_sel_o_t0;
  wire mult_sel_o_t0;
  output [1:0] multdiv_operator_o;
  wire [1:0] multdiv_operator_o;
  output [1:0] multdiv_operator_o_t0;
  wire [1:0] multdiv_operator_o_t0;
  output [1:0] multdiv_signed_mode_o;
  wire [1:0] multdiv_signed_mode_o;
  output [1:0] multdiv_signed_mode_o_t0;
  wire [1:0] multdiv_signed_mode_o_t0;
  output [4:0] rf_raddr_a_o;
  wire [4:0] rf_raddr_a_o;
  output [4:0] rf_raddr_a_o_t0;
  wire [4:0] rf_raddr_a_o_t0;
  output [4:0] rf_raddr_b_o;
  wire [4:0] rf_raddr_b_o;
  output [4:0] rf_raddr_b_o_t0;
  wire [4:0] rf_raddr_b_o_t0;
  output rf_ren_a_o;
  wire rf_ren_a_o;
  output rf_ren_a_o_t0;
  wire rf_ren_a_o_t0;
  output rf_ren_b_o;
  wire rf_ren_b_o;
  output rf_ren_b_o_t0;
  wire rf_ren_b_o_t0;
  output [4:0] rf_waddr_o;
  wire [4:0] rf_waddr_o;
  output [4:0] rf_waddr_o_t0;
  wire [4:0] rf_waddr_o_t0;
  output rf_wdata_sel_o;
  wire rf_wdata_sel_o;
  output rf_wdata_sel_o_t0;
  wire rf_wdata_sel_o_t0;
  output rf_we_o;
  wire rf_we_o;
  output rf_we_o_t0;
  wire rf_we_o_t0;
  input rst_ni;
  wire rst_ni;
  output wfi_insn_o;
  wire wfi_insn_o;
  output wfi_insn_o_t0;
  wire wfi_insn_o_t0;
  output [31:0] zimm_rs1_type_o;
  wire [31:0] zimm_rs1_type_o;
  output [31:0] zimm_rs1_type_o_t0;
  wire [31:0] zimm_rs1_type_o_t0;
  assign _0363_ = | csr_op_t0;
  assign _0365_ = | { instr_rdata_i_t0[26], instr_rdata_i_t0[13:12] };
  assign _0366_ = | instr_rdata_alu_i_t0[31:27];
  assign _0369_ = | { instr_rdata_alu_i_t0[31:25], instr_rdata_alu_i_t0[14:12] };
  assign _0371_ = | instr_rdata_alu_i_t0[6:0];
  assign _0374_ = | { instr_rdata_i_t0[31:25], instr_rdata_i_t0[14:12] };
  assign _0376_ = | instr_rdata_i_t0[31:27];
  assign _0379_ = | instr_rdata_i_t0[6:0];
  assign _0270_ = ~ csr_op_t0;
  assign _0272_ = ~ { instr_rdata_i_t0[26], instr_rdata_i_t0[13:12] };
  assign _0273_ = ~ instr_rdata_alu_i_t0[31:27];
  assign _0283_ = ~ { instr_rdata_alu_i_t0[31:25], instr_rdata_alu_i_t0[14:12] };
  assign _0288_ = ~ instr_rdata_alu_i_t0[14:12];
  assign _0293_ = ~ instr_rdata_alu_i_t0[6:0];
  assign _0297_ = ~ instr_rdata_i_t0[13:12];
  assign _0300_ = ~ instr_rdata_i_t0[31:20];
  assign _0303_ = ~ { instr_rdata_i_t0[31:25], instr_rdata_i_t0[14:12] };
  assign _0307_ = ~ instr_rdata_i_t0[31:27];
  assign _0278_ = ~ instr_rdata_i_t0[14:12];
  assign _0311_ = ~ instr_rdata_i_t0[6:0];
  assign _0682_ = csr_op & _0270_;
  assign _0686_ = { instr_rdata_i[26], instr_rdata_i[13:12] } & _0272_;
  assign _0688_ = instr_rdata_alu_i[31:27] & _0273_;
  assign _0713_ = { instr_rdata_alu_i[31:25], instr_rdata_alu_i[14:12] } & _0283_;
  assign _0743_ = instr_rdata_alu_i[14:12] & _0288_;
  assign _0763_ = instr_rdata_alu_i[6:0] & _0293_;
  assign _0800_ = instr_rdata_i[13:12] & _0297_;
  assign _0804_ = instr_rdata_i[31:20] & _0300_;
  assign _0829_ = { instr_rdata_i[31:25], instr_rdata_i[14:12] } & _0303_;
  assign _0857_ = instr_rdata_i[31:27] & _0307_;
  assign _0699_ = instr_rdata_i[14:12] & _0278_;
  assign _0874_ = instr_rdata_i[6:0] & _0311_;
  assign _0683_ = 2'h2 & _0270_;
  assign _0684_ = 2'h3 & _0270_;
  assign _0687_ = 3'h5 & _0272_;
  assign _0689_ = 5'h08 & _0273_;
  assign _0714_ = 10'h105 & _0283_;
  assign _0715_ = 10'h005 & _0283_;
  assign _0716_ = 10'h001 & _0283_;
  assign _0717_ = 10'h007 & _0283_;
  assign _0718_ = 10'h006 & _0283_;
  assign _0719_ = 10'h004 & _0283_;
  assign _0720_ = 10'h002 & _0283_;
  assign _0721_ = 10'h100 & _0283_;
  assign _0722_ = 10'h00f & _0283_;
  assign _0723_ = 10'h00e & _0283_;
  assign _0724_ = 10'h00d & _0283_;
  assign _0725_ = 10'h00c & _0283_;
  assign _0726_ = 10'h00b & _0283_;
  assign _0727_ = 10'h00a & _0283_;
  assign _0728_ = 10'h009 & _0283_;
  assign _0729_ = 10'h008 & _0283_;
  assign _0744_ = 3'h3 & _0288_;
  assign _0745_ = 3'h2 & _0288_;
  assign _0758_ = 3'h7 & _0288_;
  assign _0759_ = 3'h6 & _0288_;
  assign _0760_ = 3'h5 & _0288_;
  assign _0761_ = 3'h4 & _0288_;
  assign _0762_ = 3'h1 & _0288_;
  assign _0764_ = 7'h13 & _0293_;
  assign _0765_ = 7'h03 & _0293_;
  assign _0766_ = 7'h17 & _0293_;
  assign _0767_ = 7'h37 & _0293_;
  assign _0768_ = 7'h23 & _0293_;
  assign _0772_ = 7'h0f & _0293_;
  assign _0773_ = 7'h63 & _0293_;
  assign _0774_ = 7'h67 & _0293_;
  assign _0775_ = 7'h6f & _0293_;
  assign _0780_ = 7'h33 & _0293_;
  assign _0783_ = 7'h73 & _0293_;
  assign _0801_ = 2'h3 & _0297_;
  assign _0805_ = 12'h105 & _0300_;
  assign _0806_ = 12'h7b2 & _0300_;
  assign _0807_ = 12'h302 & _0300_;
  assign _0808_ = 12'h001 & _0300_;
  assign _0830_ = 10'h008 & _0303_;
  assign _0831_ = 10'h100 & _0303_;
  assign _0832_ = 10'h002 & _0303_;
  assign _0833_ = 10'h003 & _0303_;
  assign _0834_ = 10'h004 & _0303_;
  assign _0835_ = 10'h006 & _0303_;
  assign _0836_ = 10'h007 & _0303_;
  assign _0837_ = 10'h001 & _0303_;
  assign _0838_ = 10'h005 & _0303_;
  assign _0839_ = 10'h105 & _0303_;
  assign _0840_ = 10'h00f & _0303_;
  assign _0841_ = 10'h00e & _0303_;
  assign _0842_ = 10'h00d & _0303_;
  assign _0843_ = 10'h00c & _0303_;
  assign _0844_ = 10'h00b & _0303_;
  assign _0845_ = 10'h00a & _0303_;
  assign _0846_ = 10'h009 & _0303_;
  assign _0858_ = 5'h08 & _0307_;
  assign _0866_ = 2'h2 & _0297_;
  assign _0867_ = 2'h1 & _0297_;
  assign _0869_ = 3'h1 & _0278_;
  assign _0870_ = 3'h4 & _0278_;
  assign _0871_ = 3'h5 & _0278_;
  assign _0872_ = 3'h6 & _0278_;
  assign _0873_ = 3'h7 & _0278_;
  assign _0875_ = 7'h0f & _0311_;
  assign _0876_ = 7'h17 & _0311_;
  assign _0877_ = 7'h37 & _0311_;
  assign _0878_ = 7'h6f & _0311_;
  assign _0900_ = 7'h33 & _0311_;
  assign _0901_ = 7'h13 & _0311_;
  assign _0902_ = 7'h03 & _0311_;
  assign _0903_ = 7'h23 & _0311_;
  assign _0904_ = 7'h63 & _0311_;
  assign _0905_ = 7'h67 & _0311_;
  assign _0906_ = 7'h73 & _0311_;
  assign _1261_ = _0682_ == _0683_;
  assign _1262_ = _0682_ == _0684_;
  assign _1263_ = _0686_ == _0687_;
  assign _1264_ = _0688_ == _0689_;
  assign _1265_ = _0713_ == _0714_;
  assign _1266_ = _0713_ == _0715_;
  assign _1267_ = _0713_ == _0716_;
  assign _1268_ = _0713_ == _0717_;
  assign _1269_ = _0713_ == _0718_;
  assign _1270_ = _0713_ == _0719_;
  assign _1271_ = _0713_ == _0720_;
  assign _1272_ = _0713_ == _0721_;
  assign _1273_ = _0713_ == _0722_;
  assign _1274_ = _0713_ == _0723_;
  assign _1275_ = _0713_ == _0724_;
  assign _1276_ = _0713_ == _0725_;
  assign _1277_ = _0713_ == _0726_;
  assign _1278_ = _0713_ == _0727_;
  assign _1279_ = _0713_ == _0728_;
  assign _1280_ = _0713_ == _0729_;
  assign _1281_ = _0743_ == _0744_;
  assign _1282_ = _0743_ == _0745_;
  assign _1283_ = _0743_ == _0758_;
  assign _1284_ = _0743_ == _0759_;
  assign _1285_ = _0743_ == _0760_;
  assign _1286_ = _0743_ == _0761_;
  assign _1287_ = _0743_ == _0762_;
  assign _1288_ = _0763_ == _0764_;
  assign _1289_ = _0763_ == _0765_;
  assign _1290_ = _0763_ == _0766_;
  assign _1291_ = _0763_ == _0767_;
  assign _1292_ = _0763_ == _0768_;
  assign _1293_ = _0763_ == _0772_;
  assign _1294_ = _0763_ == _0773_;
  assign _1295_ = _0763_ == _0774_;
  assign _1296_ = _0763_ == _0775_;
  assign _1297_ = _0763_ == _0780_;
  assign _1298_ = _0763_ == _0783_;
  assign _1299_ = _0800_ == _0801_;
  assign _1300_ = _0804_ == _0805_;
  assign _1301_ = _0804_ == _0806_;
  assign _1302_ = _0804_ == _0807_;
  assign _1303_ = _0804_ == _0808_;
  assign _1304_ = _0829_ == _0830_;
  assign _1305_ = _0829_ == _0831_;
  assign _1306_ = _0829_ == _0832_;
  assign _1307_ = _0829_ == _0833_;
  assign _1308_ = _0829_ == _0834_;
  assign _1309_ = _0829_ == _0835_;
  assign _1310_ = _0829_ == _0836_;
  assign _1311_ = _0829_ == _0837_;
  assign _1312_ = _0829_ == _0838_;
  assign _1313_ = _0829_ == _0839_;
  assign _1314_ = _0829_ == _0840_;
  assign _1315_ = _0829_ == _0841_;
  assign _1316_ = _0829_ == _0842_;
  assign _1317_ = _0829_ == _0843_;
  assign _1318_ = _0829_ == _0844_;
  assign _1319_ = _0829_ == _0845_;
  assign _1320_ = _0829_ == _0846_;
  assign _1321_ = _0857_ == _0858_;
  assign _1322_ = _0800_ == _0866_;
  assign _1323_ = _0800_ == _0867_;
  assign _1324_ = _0699_ == _0869_;
  assign _1325_ = _0699_ == _0870_;
  assign _1326_ = _0699_ == _0871_;
  assign _1327_ = _0699_ == _0872_;
  assign _1328_ = _0699_ == _0873_;
  assign _1329_ = _0874_ == _0875_;
  assign _1330_ = _0874_ == _0876_;
  assign _1331_ = _0874_ == _0877_;
  assign _1332_ = _0874_ == _0878_;
  assign _1333_ = _0874_ == _0900_;
  assign _1334_ = _0874_ == _0901_;
  assign _1335_ = _0874_ == _0902_;
  assign _1336_ = _0874_ == _0903_;
  assign _1337_ = _0874_ == _0904_;
  assign _1338_ = _0874_ == _0905_;
  assign _1339_ = _0874_ == _0906_;
  assign _1444_ = _1261_ & _0363_;
  assign _1446_ = _1262_ & _0363_;
  assign _1450_ = _1263_ & _0365_;
  assign _1455_ = _1264_ & _0366_;
  assign _1490_ = _1265_ & _0369_;
  assign _1492_ = _1266_ & _0369_;
  assign _1494_ = _1267_ & _0369_;
  assign _1496_ = _1268_ & _0369_;
  assign _1498_ = _1269_ & _0369_;
  assign _1500_ = _1270_ & _0369_;
  assign _1502_ = _1271_ & _0369_;
  assign _1504_ = _1272_ & _0369_;
  assign _1474_ = _1273_ & _0369_;
  assign _1476_ = _1274_ & _0369_;
  assign _1478_ = _1275_ & _0369_;
  assign _1480_ = _1276_ & _0369_;
  assign _1482_ = _1277_ & _0369_;
  assign _1484_ = _1278_ & _0369_;
  assign _1486_ = _1279_ & _0369_;
  assign _1488_ = _1280_ & _0369_;
  assign _1520_ = _1281_ & _0370_;
  assign _1522_ = _1282_ & _0370_;
  assign _1514_ = _1283_ & _0370_;
  assign _1516_ = _1284_ & _0370_;
  assign _1510_ = _1285_ & _0370_;
  assign _1518_ = _1286_ & _0370_;
  assign _1470_ = _1287_ & _0370_;
  assign _1512_ = _1288_ & _0371_;
  assign _1534_ = _1289_ & _0371_;
  assign _1532_ = _1290_ & _0371_;
  assign _1536_ = _1291_ & _0371_;
  assign _1524_ = _1292_ & _0371_;
  assign _1472_ = _1293_ & _0371_;
  assign _1526_ = _1294_ & _0371_;
  assign _1528_ = _1295_ & _0371_;
  assign _1530_ = _1296_ & _0371_;
  assign _1508_ = _1297_ & _0371_;
  assign _1468_ = _1298_ & _0371_;
  assign _1538_ = _1299_ & _0372_;
  assign _0096_ = _1300_ & _0373_;
  assign _0079_ = _1301_ & _0373_;
  assign _0087_ = _1302_ & _0373_;
  assign _0081_ = _1303_ & _0373_;
  assign _1568_ = _1304_ & _0374_;
  assign _1570_[1] = _1305_ & _0374_;
  assign _1570_[2] = _1306_ & _0374_;
  assign _1570_[3] = _1307_ & _0374_;
  assign _1570_[4] = _1308_ & _0374_;
  assign _1570_[5] = _1309_ & _0374_;
  assign _1570_[6] = _1310_ & _0374_;
  assign _1570_[7] = _1311_ & _0374_;
  assign _1570_[8] = _1312_ & _0374_;
  assign _1570_[9] = _1313_ & _0374_;
  assign _1554_ = _1314_ & _0374_;
  assign _1556_ = _1315_ & _0374_;
  assign _1558_ = _1316_ & _0374_;
  assign _1560_ = _1317_ & _0374_;
  assign _1562_ = _1318_ & _0374_;
  assign _1564_ = _1319_ & _0374_;
  assign _1566_ = _1320_ & _0374_;
  assign _1578_[1] = _1321_ & _0376_;
  assign _1540_ = _1322_ & _0372_;
  assign _1542_ = _1323_ & _0372_;
  assign _0058_ = _1324_ & _0367_;
  assign _1582_[3] = _1325_ & _0367_;
  assign _1574_ = _1326_ & _0367_;
  assign _1582_[4] = _1327_ & _0367_;
  assign _1582_[5] = _1328_ & _0367_;
  assign _1552_ = _1329_ & _0379_;
  assign _1595_ = _1330_ & _0379_;
  assign _1597_ = _1331_ & _0379_;
  assign _1593_ = _1332_ & _0379_;
  assign _1572_ = _1333_ & _0379_;
  assign _1576_ = _1334_ & _0379_;
  assign _1584_ = _1335_ & _0379_;
  assign _0019_ = _1336_ & _0379_;
  assign _0015_ = _1337_ & _0379_;
  assign _1591_ = _1338_ & _0379_;
  assign _1544_ = _1339_ & _0379_;
  assign _0690_ = _1460_ & _1447_;
  assign _0691_ = _1448_ & _1459_;
  assign _0692_ = _1460_ & _1448_;
  assign _1141_ = _0690_ | _0691_;
  assign _1458_ = _1141_ | _0692_;
  assign _0335_ = | { _1593_, _1591_ };
  assign _0336_ = | { _1584_, _0019_ };
  assign _0337_ = | { _1530_, _1532_, _1528_ };
  assign _0338_ = | { _0058_, _0039_ };
  assign _0339_ = | { _1572_, _0019_, _0015_ };
  assign _0340_ = | { _0081_, _0087_, _0079_, _0096_, _0083_ };
  assign _0341_ = | { _1593_, _1595_, _1597_, _1576_, _1572_, _1591_ };
  assign _0342_ = | { _1554_, _1556_ };
  assign _0343_ = | { _1560_, _1558_ };
  assign _0344_ = | { _1566_, _1564_, _1562_ };
  assign _0345_ = | { _1488_, _1486_, _1484_, _1482_ };
  assign _0346_ = | { _1566_, _1560_, _1556_ };
  assign _0347_ = | { _1476_, _1480_, _1478_, _1474_ };
  assign _0348_ = | { _1506_, _1476_, _1488_, _1480_, _1478_, _1474_, _1486_, _1484_, _1482_ };
  assign _0349_ = | { _1532_, _1536_ };
  assign _0350_ = | { _1530_, _1528_ };
  assign _0351_ = | { _1584_, _1576_, _1572_, _1591_, _0019_, _0015_ };
  assign _0352_ = | { _1566_, _1560_, _1554_, _1564_, _1562_, _1558_, _1556_, _1570_, _1568_ };
  assign _0353_ = | { _1530_, _1532_, _1536_, _1528_, _1524_, _1534_ };
  assign _0354_ = | { _1542_, _1540_, _1538_ };
  assign _0355_ = | { _1586_, _1542_, _1540_ };
  assign _0356_ = | { _1586_, _1542_ };
  assign _0357_ = | { _0923_, _1496_, _1494_, _1492_ };
  assign _0358_ = | { _0927_, _1514_, _1516_ };
  assign _0359_ = | { _1510_, _1514_, _1516_ };
  assign _0360_ = | { _1512_, _1468_, _1524_, _1534_, _1508_, _1472_ };
  assign _0361_ = | { _1512_, _1508_, _1472_ };
  assign _0362_ = | { _1593_, _1595_, _1597_, _1576_, _1572_, _0943_ };
  assign _0364_ = | instr_rdata_i_t0[19:15];
  assign _0368_ = | instr_rdata_i_t0[11:7];
  assign _0370_ = | instr_rdata_alu_i_t0[14:12];
  assign _0373_ = | instr_rdata_i_t0[31:20];
  assign _0375_ = | _1578_;
  assign _0377_ = | instr_rdata_i_t0[26:25];
  assign _0372_ = | instr_rdata_i_t0[13:12];
  assign _0378_ = | { _1574_, _0058_, _0039_, _1582_[5:3] };
  assign _0367_ = | instr_rdata_i_t0[14:12];
  assign _0168_ = ~ { _1593_, _1591_ };
  assign _0169_ = ~ { _0019_, _1584_ };
  assign _0170_ = ~ { _1532_, _1530_, _1528_ };
  assign _0171_ = ~ { _0058_, _0039_ };
  assign _0172_ = ~ { _0015_, _0019_, _1572_ };
  assign _0173_ = ~ { _0081_, _0087_, _0079_, _0096_, _0083_ };
  assign _0174_ = ~ { _1597_, _1595_, _1593_, _1591_, _1576_, _1572_ };
  assign _0175_ = ~ { _1556_, _1554_ };
  assign _0176_ = ~ { _1560_, _1558_ };
  assign _0177_ = ~ { _1566_, _1564_, _1562_ };
  assign _0178_ = ~ { _1488_, _1486_, _1484_, _1482_ };
  assign _0179_ = ~ { _1566_, _1560_, _1556_ };
  assign _0180_ = ~ { _1480_, _1478_, _1476_, _1474_ };
  assign _0181_ = ~ { _1506_, _1488_, _1486_, _1484_, _1482_, _1480_, _1478_, _1476_, _1474_ };
  assign _0182_ = ~ { _1536_, _1532_ };
  assign _0183_ = ~ { _1530_, _1528_ };
  assign _0184_ = ~ { _1591_, _0015_, _0019_, _1584_, _1576_, _1572_ };
  assign _0185_ = ~ { _1570_, _1568_, _1566_, _1564_, _1562_, _1560_, _1558_, _1556_, _1554_ };
  assign _0186_ = ~ { _1536_, _1534_, _1532_, _1530_, _1528_, _1524_ };
  assign _0187_ = ~ { _1542_, _1540_, _1538_ };
  assign _0188_ = ~ { _1586_, _1542_, _1540_ };
  assign _0189_ = ~ { _1586_, _1542_ };
  assign _0211_ = ~ { _0923_, _1496_, _1494_, _1492_ };
  assign _0212_ = ~ { _1516_, _1514_, _0927_ };
  assign _0213_ = ~ { _1516_, _1514_, _1510_ };
  assign _0214_ = ~ { _1534_, _1524_, _1512_, _1508_, _1472_, _1468_ };
  assign _0215_ = ~ { _1512_, _1508_, _1472_ };
  assign _0216_ = ~ { _0943_, _1597_, _1595_, _1593_, _1576_, _1572_ };
  assign _0271_ = ~ instr_rdata_i_t0[19:15];
  assign _0279_ = ~ instr_rdata_i_t0[11:7];
  assign _0306_ = ~ _1578_;
  assign _0309_ = ~ instr_rdata_i_t0[26:25];
  assign _0310_ = ~ { _1582_[5:3], _1574_, _0058_, _0039_ };
  assign _0421_ = { _1592_, _1590_ } & _0168_;
  assign _0422_ = { _1587_, _1583_ } & _0169_;
  assign _0423_ = { _1531_, _1529_, _1527_ } & _0170_;
  assign _0424_ = { _1550_, _1451_ } & _0171_;
  assign _0425_ = { _1589_, _1587_, _1571_ } & _0172_;
  assign _0426_ = { _1549_, _1548_, _1547_, _1546_, _1545_ } & _0173_;
  assign _0427_ = { _1596_, _1594_, _1592_, _1590_, _1575_, _1571_ } & _0174_;
  assign _0428_ = { _1555_, _1553_ } & _0175_;
  assign _0429_ = { _1559_, _1557_ } & _0176_;
  assign _0430_ = { _1565_, _1563_, _1561_ } & _0177_;
  assign _0431_ = { _1487_, _1485_, _1483_, _1481_ } & _0178_;
  assign _0432_ = { _1565_, _1559_, _1555_ } & _0179_;
  assign _0433_ = { _1479_, _1477_, _1475_, _1473_ } & _0180_;
  assign _0434_ = { _1505_, _1487_, _1485_, _1483_, _1481_, _1479_, _1477_, _1475_, _1473_ } & _0181_;
  assign _0435_ = { _1535_, _1531_ } & _0182_;
  assign _0436_ = { _1529_, _1527_ } & _0183_;
  assign _0437_ = { _1590_, _1589_, _1587_, _1583_, _1575_, _1571_ } & _0184_;
  assign _0438_ = { _1569_, _1567_, _1565_, _1563_, _1561_, _1559_, _1557_, _1555_, _1553_ } & _0185_;
  assign _0439_ = { _1535_, _1533_, _1531_, _1529_, _1527_, _1523_ } & _0186_;
  assign _0440_ = { _1541_, _1539_, _1537_ } & _0187_;
  assign _0441_ = { _1585_, _1541_, _1539_ } & _0188_;
  assign _0442_ = { _1585_, _1541_ } & _0189_;
  assign _0479_ = { _0922_, _1495_, _1493_, _1491_ } & _0211_;
  assign _0480_ = { _1515_, _1513_, _0926_ } & _0212_;
  assign _0481_ = { _1515_, _1513_, _1509_ } & _0213_;
  assign _0482_ = { _1533_, _1523_, _1511_, _1507_, _1471_, _1467_ } & _0214_;
  assign _0483_ = { _1511_, _1507_, _1471_ } & _0215_;
  assign _0484_ = { _0942_, _1596_, _1594_, _1592_, _1575_, _1571_ } & _0216_;
  assign _0685_ = instr_rdata_i[19:15] & _0271_;
  assign _0700_ = instr_rdata_i[11:7] & _0279_;
  assign _0856_ = _1577_ & _0306_;
  assign _0861_ = instr_rdata_i[26:25] & _0309_;
  assign _0868_ = { _1581_[5:3], _1573_, _1550_, _1451_ } & _0310_;
  assign _0380_ = ! _0421_;
  assign _0381_ = ! _0422_;
  assign _0382_ = ! _0423_;
  assign _0383_ = ! _0424_;
  assign _0384_ = ! _0425_;
  assign _0385_ = ! _0426_;
  assign _0386_ = ! _0427_;
  assign _0387_ = ! _0428_;
  assign _0388_ = ! _0429_;
  assign _0389_ = ! _0430_;
  assign _0390_ = ! _0431_;
  assign _0391_ = ! _0432_;
  assign _0392_ = ! _0433_;
  assign _0393_ = ! _0434_;
  assign _0394_ = ! _0435_;
  assign _0395_ = ! _0436_;
  assign _0396_ = ! _0437_;
  assign _0397_ = ! _0438_;
  assign _0398_ = ! _0439_;
  assign _0399_ = ! _0440_;
  assign _0400_ = ! _0441_;
  assign _0401_ = ! _0442_;
  assign _0402_ = ! _0479_;
  assign _0403_ = ! _0480_;
  assign _0404_ = ! _0481_;
  assign _0405_ = ! _0482_;
  assign _0406_ = ! _0483_;
  assign _0407_ = ! _0484_;
  assign _0409_ = ! _0688_;
  assign _0408_ = ! _0685_;
  assign _0411_ = ! _0700_;
  assign _0412_ = ! _0713_;
  assign _0413_ = ! _0743_;
  assign _0414_ = ! _0804_;
  assign _0415_ = ! _0829_;
  assign _0416_ = ! _0856_;
  assign _0417_ = ! _0861_;
  assign _0418_ = ! _0857_;
  assign _0419_ = ! _0800_;
  assign _0420_ = ! _0868_;
  assign _0410_ = ! _0699_;
  assign _0133_ = _0380_ & _0335_;
  assign _0017_ = _0381_ & _0336_;
  assign _0136_ = _0382_ & _0337_;
  assign _0031_ = _0383_ & _0338_;
  assign rf_ren_b_o_t0 = _0384_ & _0339_;
  assign _0035_ = _0385_ & _0340_;
  assign _0142_ = _0386_ & _0341_;
  assign _0144_ = _0387_ & _0342_;
  assign _0146_ = _0388_ & _0343_;
  assign _0148_ = _0389_ & _0344_;
  assign _0089_ = _0390_ & _0345_;
  assign _0153_ = _0391_ & _0346_;
  assign _0077_ = _0392_ & _0347_;
  assign _0156_ = _0393_ & _0348_;
  assign _0158_ = _0394_ & _0349_;
  assign _0160_ = _0395_ & _0350_;
  assign _0162_ = _0396_ & _0351_;
  assign _0029_ = _0397_ & _0352_;
  assign _0167_ = _0398_ & _0353_;
  assign _0073_ = _0399_ & _0354_;
  assign _0150_ = _0400_ & _0355_;
  assign _0164_ = _0401_ & _0356_;
  assign _0324_ = _0402_ & _0357_;
  assign _0326_ = _0403_ & _0358_;
  assign _0328_ = _0404_ & _0359_;
  assign _0330_ = _0405_ & _0360_;
  assign _0332_ = _0406_ & _0361_;
  assign _0334_ = _0407_ & _0362_;
  assign _1453_ = _0409_ & _0366_;
  assign _1448_ = _0408_ & _0364_;
  assign _1466_ = _0411_ & _0368_;
  assign _1506_ = _0412_ & _0369_;
  assign _0056_ = _0413_ & _0370_;
  assign _0083_ = _0414_ & _0373_;
  assign _1570_[0] = _0415_ & _0374_;
  assign _1580_ = _0416_ & _0375_;
  assign _0914_ = _0417_ & _0377_;
  assign _1578_[0] = _0418_ & _0376_;
  assign _1586_ = _0419_ & _0372_;
  assign _0085_ = _0420_ & _0378_;
  assign _0039_ = _0410_ & _0367_;
  assign _0274_ = ~ _1443_;
  assign _0276_ = ~ _1464_;
  assign _0275_ = ~ _1445_;
  assign _0277_ = ~ _1465_;
  assign _0693_ = _1444_ & _0275_;
  assign _0696_ = _1448_ & _0277_;
  assign _0694_ = _1446_ & _0274_;
  assign _0697_ = _1466_ & _0276_;
  assign _0695_ = _1444_ & _1446_;
  assign _0698_ = _1448_ & _1466_;
  assign _1142_ = _0693_ | _0694_;
  assign _1143_ = _0696_ | _0697_;
  assign _1460_ = _1142_ | _0695_;
  assign _1462_ = _1143_ | _0698_;
  assign _0217_ = ~ { _0155_, _0155_, _0155_, _0155_, _0155_, _0155_ };
  assign _0218_ = ~ { _1493_, _1493_, _1493_, _1493_, _1493_, _1493_ };
  assign _0219_ = ~ { _1491_, _1491_, _1491_, _1491_, _1491_, _1491_ };
  assign _0220_ = ~ { _0922_, _0922_, _0922_, _0922_, _0922_, _0922_ };
  assign _0221_ = ~ { _1497_, _1497_, _1497_, _1497_, _1497_, _1497_ };
  assign _0222_ = ~ { _1503_, _1503_, _1503_, _1503_, _1503_, _1503_ };
  assign _0223_ = ~ { _1501_, _1501_, _1501_, _1501_, _1501_, _1501_ };
  assign _0224_ = ~ { _0924_, _0924_, _0924_, _0924_, _0924_, _0924_ };
  assign _0225_ = ~ { _0323_, _0323_, _0323_, _0323_, _0323_, _0323_ };
  assign _0226_ = ~ { _1509_, _1509_, _1509_, _1509_, _1509_, _1509_ };
  assign _0228_ = ~ { _0926_, _0926_, _0926_, _0926_, _0926_, _0926_ };
  assign _0230_ = ~ { _1521_, _1521_, _1521_, _1521_, _1521_, _1521_ };
  assign _0231_ = ~ { _0928_, _0928_, _0928_, _0928_, _0928_, _0928_ };
  assign _0232_ = ~ { _0325_, _0325_, _0325_, _0325_, _0325_, _0325_ };
  assign _0233_ = ~ { _1515_, _1515_, _1515_, _1515_, _1515_, _1515_ };
  assign _0227_ = ~ { _1513_, _1513_, _1513_, _1513_, _1513_, _1513_ };
  assign _0229_ = ~ { _1517_, _1517_, _1517_, _1517_, _1517_, _1517_ };
  assign _0235_ = ~ { _0930_, _0930_, _0930_, _0930_, _0930_, _0930_ };
  assign _0236_ = ~ { _0327_, _0327_, _0327_, _0327_, _0327_, _0327_ };
  assign _0201_ = ~ _1525_;
  assign _0237_ = ~ _0932_;
  assign _0238_ = ~ { _1471_, _1471_ };
  assign _0239_ = ~ { _1467_, _1467_ };
  assign _0240_ = ~ { _1525_, _1525_ };
  assign _0241_ = ~ { _0135_, _0135_ };
  assign _0242_ = ~ { _0329_, _0329_ };
  assign _0243_ = ~ { _1507_, _1507_, _1507_, _1507_, _1507_, _1507_ };
  assign _0244_ = ~ { _1471_, _1471_, _1471_, _1471_, _1471_, _1471_ };
  assign _0245_ = ~ { _1525_, _1525_, _1525_, _1525_, _1525_, _1525_ };
  assign _0246_ = ~ { _0166_, _0166_, _0166_, _0166_, _0166_, _0166_ };
  assign _0247_ = ~ { _0331_, _0331_, _0331_, _0331_, _0331_, _0331_ };
  assign _0248_ = ~ { _0157_, _0157_, _0157_ };
  assign _0249_ = ~ { _0159_, _0159_, _0159_ };
  assign _0250_ = ~ { _1525_, _1525_, _1525_ };
  assign _0251_ = ~ { _0934_, _0934_, _0934_ };
  assign _0252_ = ~ { _1471_, _1471_, _1471_ };
  assign _0253_ = ~ { _1529_, _1529_, _1529_ };
  assign _0254_ = ~ { _0936_, _0936_, _0936_ };
  assign _0255_ = ~ { _1537_, _1537_ };
  assign _0257_ = ~ { _0938_, _0938_ };
  assign _0258_ = ~ { _1563_, _1563_ };
  assign _0259_ = ~ { _0152_, _0152_ };
  assign _0260_ = ~ { _0143_, _0143_ };
  assign _0261_ = ~ { _0147_, _0147_ };
  assign _0262_ = ~ { _0940_, _0940_ };
  assign _0263_ = ~ _1573_;
  assign _0203_ = ~ _1539_;
  assign _0264_ = ~ { _1585_, _1585_ };
  assign _0256_ = ~ { _1541_, _1541_ };
  assign _0265_ = ~ _1571_;
  assign _0266_ = ~ _0942_;
  assign _0268_ = ~ _0944_;
  assign _0269_ = ~ _0333_;
  assign _0280_ = ~ { instr_rdata_alu_i[14], instr_rdata_alu_i[14] };
  assign _0281_ = ~ { _1456_, _1456_ };
  assign _0234_ = ~ { _1456_, _1456_, _1456_, _1456_, _1456_, _1456_ };
  assign _0282_ = ~ { _1469_, _1469_, _1469_ };
  assign _0284_ = ~ instr_rdata_alu_i[26];
  assign _0285_ = ~ { instr_rdata_alu_i[26], instr_rdata_alu_i[26], instr_rdata_alu_i[26], instr_rdata_alu_i[26], instr_rdata_alu_i[26], instr_rdata_alu_i[26] };
  assign _0286_ = ~ { _1454_, _1454_, _1454_, _1454_, _1454_, _1454_ };
  assign _0287_ = ~ { _1452_, _1452_, _1452_, _1452_, _1452_, _1452_ };
  assign _0289_ = ~ { instr_rdata_alu_i[14], instr_rdata_alu_i[14], instr_rdata_alu_i[14] };
  assign _0290_ = ~ { instr_first_cycle_i, instr_first_cycle_i };
  assign _0291_ = ~ { instr_first_cycle_i, instr_first_cycle_i, instr_first_cycle_i, instr_first_cycle_i, instr_first_cycle_i, instr_first_cycle_i };
  assign _0292_ = ~ { instr_first_cycle_i, instr_first_cycle_i, instr_first_cycle_i };
  assign _0294_ = ~ { _1527_, _1527_ };
  assign _0199_ = ~ _1507_;
  assign _0296_ = ~ illegal_c_insn_i;
  assign _0299_ = ~ _1461_;
  assign _0301_ = ~ _1451_;
  assign _0302_ = ~ { _1451_, _1451_ };
  assign _0304_ = ~ _1449_;
  assign _0305_ = ~ { _1449_, _1449_ };
  assign _0308_ = ~ instr_rdata_i[26];
  assign _0298_ = ~ instr_rdata_i[14];
  assign _0267_ = ~ _1589_;
  assign _0210_ = ~ _1583_;
  assign _0312_ = ~ { _0134_, _0134_ };
  assign _0313_ = ~ { _1571_, _1571_ };
  assign _0208_ = ~ _1543_;
  assign _0207_ = ~ _1551_;
  assign _0314_ = ~ { _1543_, _1543_ };
  assign _0209_ = ~ _1587_;
  assign _0315_ = ~ { _1457_, _1457_ };
  assign _0316_ = ~ { branch_taken_i, branch_taken_i, branch_taken_i };
  assign _0295_ = ~ illegal_insn_o;
  assign _0958_ = { _0156_, _0156_, _0156_, _0156_, _0156_, _0156_ } | _0217_;
  assign _0961_ = { _1494_, _1494_, _1494_, _1494_, _1494_, _1494_ } | _0218_;
  assign _0964_ = { _1492_, _1492_, _1492_, _1492_, _1492_, _1492_ } | _0219_;
  assign _0967_ = { _0923_, _0923_, _0923_, _0923_, _0923_, _0923_ } | _0220_;
  assign _0970_ = { _1498_, _1498_, _1498_, _1498_, _1498_, _1498_ } | _0221_;
  assign _0973_ = { _1504_, _1504_, _1504_, _1504_, _1504_, _1504_ } | _0222_;
  assign _0976_ = { _1502_, _1502_, _1502_, _1502_, _1502_, _1502_ } | _0223_;
  assign _0979_ = { _0925_, _0925_, _0925_, _0925_, _0925_, _0925_ } | _0224_;
  assign _0982_ = { _0324_, _0324_, _0324_, _0324_, _0324_, _0324_ } | _0225_;
  assign _0985_ = { _1510_, _1510_, _1510_, _1510_, _1510_, _1510_ } | _0226_;
  assign _0991_ = { _0927_, _0927_, _0927_, _0927_, _0927_, _0927_ } | _0228_;
  assign _0997_ = { _1522_, _1522_, _1522_, _1522_, _1522_, _1522_ } | _0230_;
  assign _1000_ = { _0929_, _0929_, _0929_, _0929_, _0929_, _0929_ } | _0231_;
  assign _1003_ = { _0326_, _0326_, _0326_, _0326_, _0326_, _0326_ } | _0232_;
  assign _1006_ = { _1516_, _1516_, _1516_, _1516_, _1516_, _1516_ } | _0233_;
  assign _0988_ = { _1514_, _1514_, _1514_, _1514_, _1514_, _1514_ } | _0227_;
  assign _0994_ = { _1518_, _1518_, _1518_, _1518_, _1518_, _1518_ } | _0229_;
  assign _1013_ = { _0931_, _0931_, _0931_, _0931_, _0931_, _0931_ } | _0235_;
  assign _1016_ = { _0328_, _0328_, _0328_, _0328_, _0328_, _0328_ } | _0236_;
  assign _1022_ = _0933_ | _0237_;
  assign _1025_ = { _1472_, _1472_ } | _0238_;
  assign _1028_ = { _1468_, _1468_ } | _0239_;
  assign _1031_ = { _1526_, _1526_ } | _0240_;
  assign _1034_ = { _0136_, _0136_ } | _0241_;
  assign _1037_ = { _0330_, _0330_ } | _0242_;
  assign _1040_ = { _1508_, _1508_, _1508_, _1508_, _1508_, _1508_ } | _0243_;
  assign _1043_ = { _1472_, _1472_, _1472_, _1472_, _1472_, _1472_ } | _0244_;
  assign _1046_ = { _1526_, _1526_, _1526_, _1526_, _1526_, _1526_ } | _0245_;
  assign _1049_ = { _0167_, _0167_, _0167_, _0167_, _0167_, _0167_ } | _0246_;
  assign _1052_ = { _0332_, _0332_, _0332_, _0332_, _0332_, _0332_ } | _0247_;
  assign _1055_ = { _0158_, _0158_, _0158_ } | _0248_;
  assign _1058_ = { _0160_, _0160_, _0160_ } | _0249_;
  assign _1061_ = { _1526_, _1526_, _1526_ } | _0250_;
  assign _1064_ = { _0935_, _0935_, _0935_ } | _0251_;
  assign _1067_ = { _1472_, _1472_, _1472_ } | _0252_;
  assign _1070_ = { _1530_, _1530_, _1530_ } | _0253_;
  assign _1073_ = { _0937_, _0937_, _0937_ } | _0254_;
  assign _1076_ = { _1538_, _1538_ } | _0255_;
  assign _1082_ = { _0939_, _0939_ } | _0257_;
  assign _1085_ = { _1564_, _1564_ } | _0258_;
  assign _1088_ = { _0153_, _0153_ } | _0259_;
  assign _1091_ = { _0144_, _0144_ } | _0260_;
  assign _1094_ = { _0148_, _0148_ } | _0261_;
  assign _1097_ = { _0941_, _0941_ } | _0262_;
  assign _1101_ = _1574_ | _0263_;
  assign _1104_ = _1540_ | _0203_;
  assign _1107_ = { _1586_, _1586_ } | _0264_;
  assign _1079_ = { _1542_, _1542_ } | _0256_;
  assign _1115_ = _1552_ | _0207_;
  assign _1121_ = _1572_ | _0265_;
  assign _1124_ = _0943_ | _0266_;
  assign _1134_ = _0945_ | _0268_;
  assign _1137_ = _0334_ | _0269_;
  assign _1111_ = _1544_ | _0208_;
  assign _1144_ = { instr_rdata_alu_i_t0[14], instr_rdata_alu_i_t0[14] } | _0280_;
  assign _1147_ = { _0056_, _0056_ } | _0281_;
  assign _1010_ = { _0056_, _0056_, _0056_, _0056_, _0056_, _0056_ } | _0234_;
  assign _1151_ = { _1470_, _1470_, _1470_ } | _0282_;
  assign _1154_ = instr_rdata_alu_i_t0[26] | _0284_;
  assign _1155_ = { instr_rdata_alu_i_t0[26], instr_rdata_alu_i_t0[26], instr_rdata_alu_i_t0[26], instr_rdata_alu_i_t0[26], instr_rdata_alu_i_t0[26], instr_rdata_alu_i_t0[26] } | _0285_;
  assign _1158_ = { _1455_, _1455_, _1455_, _1455_, _1455_, _1455_ } | _0286_;
  assign _1161_ = { _1453_, _1453_, _1453_, _1453_, _1453_, _1453_ } | _0287_;
  assign _1164_ = { instr_rdata_alu_i_t0[14], instr_rdata_alu_i_t0[14], instr_rdata_alu_i_t0[14] } | _0289_;
  assign _1167_ = { instr_first_cycle_i_t0, instr_first_cycle_i_t0 } | _0290_;
  assign _1170_ = { instr_first_cycle_i_t0, instr_first_cycle_i_t0, instr_first_cycle_i_t0, instr_first_cycle_i_t0, instr_first_cycle_i_t0, instr_first_cycle_i_t0 } | _0291_;
  assign _1173_ = { instr_first_cycle_i_t0, instr_first_cycle_i_t0, instr_first_cycle_i_t0 } | _0292_;
  assign _1176_ = { _1528_, _1528_ } | _0294_;
  assign _1019_ = _1508_ | _0199_;
  assign _1181_ = illegal_c_insn_i_t0 | _0296_;
  assign _1182_ = _1462_ | _0299_;
  assign _1183_ = _0039_ | _0301_;
  assign _1186_ = { _0039_, _0039_ } | _0302_;
  assign _1189_ = _1450_ | _0304_;
  assign _1190_ = { _1450_, _1450_ } | _0305_;
  assign _1195_ = instr_rdata_i_t0[26] | _0308_;
  assign _1131_ = _0015_ | _0267_;
  assign _1127_ = _1584_ | _0210_;
  assign _1198_ = { _0017_, _0017_ } | _0312_;
  assign _1201_ = { _1572_, _1572_ } | _0313_;
  assign _1205_ = { _1544_, _1544_ } | _0314_;
  assign _1208_ = { _1458_, _1458_ } | _0315_;
  assign _1211_ = { branch_taken_i_t0, branch_taken_i_t0, branch_taken_i_t0 } | _0316_;
  assign _1180_ = illegal_insn_o_t0 | _0295_;
  assign _0959_ = { _0156_, _0156_, _0156_, _0156_, _0156_, _0156_ } | { _0155_, _0155_, _0155_, _0155_, _0155_, _0155_ };
  assign _0962_ = { _1494_, _1494_, _1494_, _1494_, _1494_, _1494_ } | { _1493_, _1493_, _1493_, _1493_, _1493_, _1493_ };
  assign _0965_ = { _1492_, _1492_, _1492_, _1492_, _1492_, _1492_ } | { _1491_, _1491_, _1491_, _1491_, _1491_, _1491_ };
  assign _0968_ = { _0923_, _0923_, _0923_, _0923_, _0923_, _0923_ } | { _0922_, _0922_, _0922_, _0922_, _0922_, _0922_ };
  assign _0971_ = { _1498_, _1498_, _1498_, _1498_, _1498_, _1498_ } | { _1497_, _1497_, _1497_, _1497_, _1497_, _1497_ };
  assign _0974_ = { _1504_, _1504_, _1504_, _1504_, _1504_, _1504_ } | { _1503_, _1503_, _1503_, _1503_, _1503_, _1503_ };
  assign _0977_ = { _1502_, _1502_, _1502_, _1502_, _1502_, _1502_ } | { _1501_, _1501_, _1501_, _1501_, _1501_, _1501_ };
  assign _0980_ = { _0925_, _0925_, _0925_, _0925_, _0925_, _0925_ } | { _0924_, _0924_, _0924_, _0924_, _0924_, _0924_ };
  assign _0983_ = { _0324_, _0324_, _0324_, _0324_, _0324_, _0324_ } | { _0323_, _0323_, _0323_, _0323_, _0323_, _0323_ };
  assign _0986_ = { _1510_, _1510_, _1510_, _1510_, _1510_, _1510_ } | { _1509_, _1509_, _1509_, _1509_, _1509_, _1509_ };
  assign _0992_ = { _0927_, _0927_, _0927_, _0927_, _0927_, _0927_ } | { _0926_, _0926_, _0926_, _0926_, _0926_, _0926_ };
  assign _0998_ = { _1522_, _1522_, _1522_, _1522_, _1522_, _1522_ } | { _1521_, _1521_, _1521_, _1521_, _1521_, _1521_ };
  assign _1001_ = { _0929_, _0929_, _0929_, _0929_, _0929_, _0929_ } | { _0928_, _0928_, _0928_, _0928_, _0928_, _0928_ };
  assign _1004_ = { _0326_, _0326_, _0326_, _0326_, _0326_, _0326_ } | { _0325_, _0325_, _0325_, _0325_, _0325_, _0325_ };
  assign _1007_ = { _1516_, _1516_, _1516_, _1516_, _1516_, _1516_ } | { _1515_, _1515_, _1515_, _1515_, _1515_, _1515_ };
  assign _0989_ = { _1514_, _1514_, _1514_, _1514_, _1514_, _1514_ } | { _1513_, _1513_, _1513_, _1513_, _1513_, _1513_ };
  assign _0995_ = { _1518_, _1518_, _1518_, _1518_, _1518_, _1518_ } | { _1517_, _1517_, _1517_, _1517_, _1517_, _1517_ };
  assign _1014_ = { _0931_, _0931_, _0931_, _0931_, _0931_, _0931_ } | { _0930_, _0930_, _0930_, _0930_, _0930_, _0930_ };
  assign _1017_ = { _0328_, _0328_, _0328_, _0328_, _0328_, _0328_ } | { _0327_, _0327_, _0327_, _0327_, _0327_, _0327_ };
  assign _1021_ = _1526_ | _1525_;
  assign _1023_ = _0933_ | _0932_;
  assign _1026_ = { _1472_, _1472_ } | { _1471_, _1471_ };
  assign _1029_ = { _1468_, _1468_ } | { _1467_, _1467_ };
  assign _1032_ = { _1526_, _1526_ } | { _1525_, _1525_ };
  assign _1035_ = { _0136_, _0136_ } | { _0135_, _0135_ };
  assign _1038_ = { _0330_, _0330_ } | { _0329_, _0329_ };
  assign _1041_ = { _1508_, _1508_, _1508_, _1508_, _1508_, _1508_ } | { _1507_, _1507_, _1507_, _1507_, _1507_, _1507_ };
  assign _1044_ = { _1472_, _1472_, _1472_, _1472_, _1472_, _1472_ } | { _1471_, _1471_, _1471_, _1471_, _1471_, _1471_ };
  assign _1047_ = { _1526_, _1526_, _1526_, _1526_, _1526_, _1526_ } | { _1525_, _1525_, _1525_, _1525_, _1525_, _1525_ };
  assign _1050_ = { _0167_, _0167_, _0167_, _0167_, _0167_, _0167_ } | { _0166_, _0166_, _0166_, _0166_, _0166_, _0166_ };
  assign _1053_ = { _0332_, _0332_, _0332_, _0332_, _0332_, _0332_ } | { _0331_, _0331_, _0331_, _0331_, _0331_, _0331_ };
  assign _1056_ = { _0158_, _0158_, _0158_ } | { _0157_, _0157_, _0157_ };
  assign _1059_ = { _0160_, _0160_, _0160_ } | { _0159_, _0159_, _0159_ };
  assign _1062_ = { _1526_, _1526_, _1526_ } | { _1525_, _1525_, _1525_ };
  assign _1065_ = { _0935_, _0935_, _0935_ } | { _0934_, _0934_, _0934_ };
  assign _1068_ = { _1472_, _1472_, _1472_ } | { _1471_, _1471_, _1471_ };
  assign _1071_ = { _1530_, _1530_, _1530_ } | { _1529_, _1529_, _1529_ };
  assign _1074_ = { _0937_, _0937_, _0937_ } | { _0936_, _0936_, _0936_ };
  assign _1077_ = { _1538_, _1538_ } | { _1537_, _1537_ };
  assign _1083_ = { _0939_, _0939_ } | { _0938_, _0938_ };
  assign _1086_ = { _1564_, _1564_ } | { _1563_, _1563_ };
  assign _1089_ = { _0153_, _0153_ } | { _0152_, _0152_ };
  assign _1092_ = { _0144_, _0144_ } | { _0143_, _0143_ };
  assign _1095_ = { _0148_, _0148_ } | { _0147_, _0147_ };
  assign _1098_ = { _0941_, _0941_ } | { _0940_, _0940_ };
  assign _1102_ = _1574_ | _1573_;
  assign _1105_ = _1540_ | _1539_;
  assign _1108_ = { _1586_, _1586_ } | { _1585_, _1585_ };
  assign _1080_ = { _1542_, _1542_ } | { _1541_, _1541_ };
  assign _1114_ = _0133_ | _0132_;
  assign _1116_ = _1552_ | _1551_;
  assign _1120_ = _1576_ | _1575_;
  assign _1122_ = _1572_ | _1571_;
  assign _1125_ = _0943_ | _0942_;
  assign _1130_ = _1591_ | _1590_;
  assign _1135_ = _0945_ | _0944_;
  assign _1138_ = _0334_ | _0333_;
  assign _1145_ = { instr_rdata_alu_i_t0[14], instr_rdata_alu_i_t0[14] } | { instr_rdata_alu_i[14], instr_rdata_alu_i[14] };
  assign _1148_ = { _0056_, _0056_ } | { _1456_, _1456_ };
  assign _1011_ = { _0056_, _0056_, _0056_, _0056_, _0056_, _0056_ } | { _1456_, _1456_, _1456_, _1456_, _1456_, _1456_ };
  assign _1152_ = { _1470_, _1470_, _1470_ } | { _1469_, _1469_, _1469_ };
  assign _1156_ = { instr_rdata_alu_i_t0[26], instr_rdata_alu_i_t0[26], instr_rdata_alu_i_t0[26], instr_rdata_alu_i_t0[26], instr_rdata_alu_i_t0[26], instr_rdata_alu_i_t0[26] } | { instr_rdata_alu_i[26], instr_rdata_alu_i[26], instr_rdata_alu_i[26], instr_rdata_alu_i[26], instr_rdata_alu_i[26], instr_rdata_alu_i[26] };
  assign _1159_ = { _1455_, _1455_, _1455_, _1455_, _1455_, _1455_ } | { _1454_, _1454_, _1454_, _1454_, _1454_, _1454_ };
  assign _1162_ = { _1453_, _1453_, _1453_, _1453_, _1453_, _1453_ } | { _1452_, _1452_, _1452_, _1452_, _1452_, _1452_ };
  assign _1165_ = { instr_rdata_alu_i_t0[14], instr_rdata_alu_i_t0[14], instr_rdata_alu_i_t0[14] } | { instr_rdata_alu_i[14], instr_rdata_alu_i[14], instr_rdata_alu_i[14] };
  assign _1168_ = { instr_first_cycle_i_t0, instr_first_cycle_i_t0 } | { instr_first_cycle_i, instr_first_cycle_i };
  assign _1171_ = { instr_first_cycle_i_t0, instr_first_cycle_i_t0, instr_first_cycle_i_t0, instr_first_cycle_i_t0, instr_first_cycle_i_t0, instr_first_cycle_i_t0 } | { instr_first_cycle_i, instr_first_cycle_i, instr_first_cycle_i, instr_first_cycle_i, instr_first_cycle_i, instr_first_cycle_i };
  assign _1174_ = { instr_first_cycle_i_t0, instr_first_cycle_i_t0, instr_first_cycle_i_t0 } | { instr_first_cycle_i, instr_first_cycle_i, instr_first_cycle_i };
  assign _1177_ = { _1528_, _1528_ } | { _1527_, _1527_ };
  assign _1020_ = _1508_ | _1507_;
  assign _1179_ = _1468_ | _1467_;
  assign _1184_ = _0039_ | _1451_;
  assign _1187_ = { _0039_, _0039_ } | { _1451_, _1451_ };
  assign _1100_ = _0058_ | _1550_;
  assign _1191_ = { _1450_, _1450_ } | { _1449_, _1449_ };
  assign _1194_ = _1580_ | _1579_;
  assign _1196_ = _1578_[0] | _1577_[0];
  assign _1197_ = _0150_ | _0149_;
  assign _1132_ = _0015_ | _1589_;
  assign _1128_ = _1584_ | _1583_;
  assign _1199_ = { _0017_, _0017_ } | { _0134_, _0134_ };
  assign _1202_ = { _1572_, _1572_ } | { _1571_, _1571_ };
  assign _1112_ = _1544_ | _1543_;
  assign _1206_ = { _1544_, _1544_ } | { _1543_, _1543_ };
  assign _1209_ = { _1458_, _1458_ } | { _1457_, _1457_ };
  assign _1212_ = { branch_taken_i_t0, branch_taken_i_t0, branch_taken_i_t0 } | { branch_taken_i, branch_taken_i, branch_taken_i };
  assign _0485_ = 6'h00 & _0958_;
  assign _0488_ = 6'h00 & _0961_;
  assign _0491_ = _1343_ & _0964_;
  assign _0494_ = _1345_ & _0967_;
  assign _0497_ = 6'h00 & _0970_;
  assign _0500_ = 6'h00 & _0973_;
  assign _0503_ = _1351_ & _0976_;
  assign _0506_ = _1353_ & _0979_;
  assign _0509_ = _1355_ & _0982_;
  assign _0512_ = 6'h00 & _0985_;
  assign _0515_ = 6'h00 & _0988_;
  assign _0518_ = _1359_ & _0991_;
  assign _0524_ = 6'h00 & _0997_;
  assign _0527_ = _1365_ & _1000_;
  assign _0530_ = _1367_ & _1003_;
  assign _0533_ = 6'h00 & _1006_;
  assign _0536_ = _1369_ & _0988_;
  assign _0521_ = 6'h00 & _0994_;
  assign _0542_ = _1375_ & _1013_;
  assign _0545_ = _1377_ & _1016_;
  assign _0548_ = instr_rdata_alu_i_t0[14] & _1019_;
  assign _0552_ = _1381_ & _1022_;
  assign _0555_ = 2'h0 & _1025_;
  assign _0558_ = _1383_ & _1028_;
  assign _0561_ = 2'h0 & _1031_;
  assign _0564_ = _1387_ & _1034_;
  assign _0567_ = _1389_ & _1037_;
  assign _0570_ = _0121_ & _1040_;
  assign _0573_ = _1391_ & _1043_;
  assign _0576_ = 6'h00 & _1046_;
  assign _0579_ = _1394_ & _1049_;
  assign _0582_ = _1396_ & _1052_;
  assign _0585_ = _0117_ & _1055_;
  assign _0588_ = 3'h0 & _1058_;
  assign _0591_ = _1400_ & _1061_;
  assign _0594_ = _1402_ & _1064_;
  assign _0597_ = _0103_ & _1067_;
  assign _0600_ = 3'h0 & _1070_;
  assign _0603_ = _1406_ & _1073_;
  assign _0606_ = 2'h0 & _1076_;
  assign _0609_ = 2'h0 & _1079_;
  assign _0612_ = _1410_ & _1082_;
  assign _0615_ = 2'h0 & _1085_;
  assign _0618_ = _1412_ & _1088_;
  assign _0621_ = 2'h0 & _1091_;
  assign _0624_ = 2'h0 & _1094_;
  assign _0627_ = _1416_ & _1097_;
  assign _0632_ = _1418_ & _1101_;
  assign _0635_ = _0164_ & _1104_;
  assign _0638_ = 2'h0 & _1107_;
  assign _0641_ = _1421_ & _1079_;
  assign _0643_ = _0142_ & _1111_;
  assign _0648_ = _1424_ & _1115_;
  assign _0651_ = _0133_ & _1115_;
  assign _0654_ = _0031_ & _1111_;
  assign _0659_ = _1429_ & _1121_;
  assign _0662_ = _1431_ & _1124_;
  assign _0665_ = _0115_ & _1127_;
  assign _0670_ = _1437_ & _1131_;
  assign _0673_ = _1439_ & _1134_;
  assign _0676_ = _1441_ & _1137_;
  assign _0679_ = _0162_ & _1111_;
  assign _0701_ = 2'h0 & _1144_;
  assign _0704_ = _0125_ & _1147_;
  assign _0707_ = 2'h0 & _1147_;
  assign _0539_ = 6'h00 & _1010_;
  assign _0710_ = 3'h0 & _1151_;
  assign _0730_ = _0077_ & _1154_;
  assign _0732_ = _0089_ & _1154_;
  assign _0734_ = _0005_ & _1155_;
  assign _0737_ = 6'h00 & _1158_;
  assign _0740_ = _0001_ & _1161_;
  assign _0746_ = 3'h0 & _1164_;
  assign _0749_ = 2'h0 & _1167_;
  assign _0752_ = 6'h00 & _1170_;
  assign _0755_ = _0103_ & _1173_;
  assign _0769_ = 2'h0 & _1176_;
  assign _0784_ = rf_wdata_sel_o_t0 & _1180_;
  assign _0786_ = _0015_ & _1180_;
  assign _0788_ = _0025_ & _1180_;
  assign _0790_ = _0023_ & _1180_;
  assign _0792_ = _0019_ & _1180_;
  assign _0794_ = _0017_ & _1180_;
  assign _0796_ = _0027_ & _1180_;
  assign _0798_ = _0021_ & _1181_;
  assign _0802_ = _0035_ & _1182_;
  assign _0809_ = _0073_ & _1183_;
  assign _0822_ = instr_rdata_i_t0[14] & _1183_;
  assign _0824_ = _0075_ & _1186_;
  assign _0847_ = _0029_ & _1189_;
  assign _0849_ = _0093_ & _1190_;
  assign _0852_ = _0091_ & _1190_;
  assign _0859_ = _0011_ & _1195_;
  assign _0881_ = 2'h0 & _1198_;
  assign _0884_ = 2'h0 & _1201_;
  assign _0908_ = 2'h0 & _1205_;
  assign _0911_ = csr_op_t0 & _1208_;
  assign _0915_ = 3'h0 & _1211_;
  assign _0918_ = mult_sel_o_t0 & _1180_;
  assign _0920_ = div_sel_o_t0 & _1180_;
  assign _0486_ = 6'h00 & _0959_;
  assign _0489_ = 6'h00 & _0962_;
  assign _0492_ = 6'h00 & _0965_;
  assign _0495_ = _1341_ & _0968_;
  assign _0498_ = 6'h00 & _0971_;
  assign _0501_ = 6'h00 & _0974_;
  assign _0504_ = 6'h00 & _0977_;
  assign _0507_ = _1349_ & _0980_;
  assign _0510_ = _1347_ & _0983_;
  assign _0513_ = _0127_ & _0986_;
  assign _0519_ = _1357_ & _0992_;
  assign _0525_ = 6'h00 & _0998_;
  assign _0528_ = _1363_ & _1001_;
  assign _0531_ = _1361_ & _1004_;
  assign _0534_ = 6'h00 & _1007_;
  assign _0516_ = 6'h00 & _0989_;
  assign _0522_ = 6'h00 & _0995_;
  assign _0543_ = _1373_ & _1014_;
  assign _0546_ = _1371_ & _1017_;
  assign _0550_ = instr_first_cycle_i_t0 & _1021_;
  assign _0553_ = _1379_ & _1023_;
  assign _0556_ = _0108_ & _1026_;
  assign _0559_ = _0119_ & _1029_;
  assign _0562_ = _0098_ & _1032_;
  assign _0565_ = 2'h0 & _1035_;
  assign _0568_ = _1385_ & _1038_;
  assign _0571_ = _0003_ & _1041_;
  assign _0574_ = _0009_ & _1044_;
  assign _0577_ = _0111_ & _1047_;
  assign _0580_ = 6'h00 & _1050_;
  assign _0583_ = _1393_ & _1053_;
  assign _0586_ = 3'h0 & _1056_;
  assign _0589_ = 3'h0 & _1059_;
  assign _0592_ = _0106_ & _1062_;
  assign _0595_ = _1398_ & _1065_;
  assign _0598_ = _0113_ & _1068_;
  assign _0601_ = 3'h0 & _1071_;
  assign _0604_ = _1404_ & _1074_;
  assign _0607_ = 2'h0 & _1077_;
  assign _0613_ = _1408_ & _1083_;
  assign _0616_ = 2'h0 & _1086_;
  assign _0619_ = 2'h0 & _1089_;
  assign _0622_ = 2'h0 & _1092_;
  assign _0625_ = 2'h0 & _1095_;
  assign _0628_ = _1414_ & _1098_;
  assign _0630_ = _0131_ & _1100_;
  assign _0633_ = _0007_ & _1102_;
  assign _0636_ = instr_rdata_i_t0[14] & _1105_;
  assign _0639_ = 2'h0 & _1108_;
  assign _0610_ = 2'h0 & _1080_;
  assign _0644_ = _0039_ & _1112_;
  assign _0646_ = instr_first_cycle_i_t0 & _1114_;
  assign _0652_ = _0058_ & _1116_;
  assign _0655_ = _0033_ & _1112_;
  assign _0657_ = _0129_ & _1120_;
  assign _0660_ = _0013_ & _1122_;
  assign _0663_ = _1427_ & _1125_;
  assign _0666_ = _0123_ & _1128_;
  assign _0668_ = _0039_ & _1130_;
  assign _0671_ = _0085_ & _1132_;
  assign _0674_ = _1435_ & _1135_;
  assign _0677_ = _1433_ & _1138_;
  assign _0680_ = _0069_ & _1112_;
  assign _0702_ = 2'h0 & _1145_;
  assign _0705_ = 2'h0 & _1148_;
  assign _0540_ = 6'h00 & _1011_;
  assign _0711_ = 3'h0 & _1152_;
  assign _0735_ = 6'h00 & _1156_;
  assign _0738_ = 6'h00 & _1159_;
  assign _0741_ = 6'h00 & _1162_;
  assign _0747_ = 3'h0 & _1165_;
  assign _0750_ = 2'h0 & _1168_;
  assign _0753_ = _0101_ & _1171_;
  assign _0756_ = 3'h0 & _1174_;
  assign _0770_ = 2'h0 & _1177_;
  assign _0776_ = _0045_ & _1020_;
  assign _0778_ = _0063_ & _1020_;
  assign _0781_ = _0056_ & _1179_;
  assign _0810_ = _0037_ & _1184_;
  assign _0812_ = _0096_ & _1184_;
  assign _0814_ = _0083_ & _1184_;
  assign _0816_ = _0079_ & _1184_;
  assign _0818_ = _0087_ & _1184_;
  assign _0820_ = _0081_ & _1184_;
  assign _0825_ = 2'h0 & _1187_;
  assign _0827_ = instr_first_cycle_i_t0 & _1100_;
  assign _0850_ = 2'h0 & _1191_;
  assign _0854_ = _0914_ & _1194_;
  assign _0862_ = _0914_ & _1196_;
  assign _0864_ = instr_rdata_i_t0[14] & _1197_;
  assign _0879_ = instr_rdata_i_t0[14] & _1128_;
  assign _0882_ = _0043_ & _1199_;
  assign _0885_ = _0067_ & _1202_;
  assign _0887_ = _0065_ & _1202_;
  assign _0890_ = _0071_ & _1112_;
  assign _0892_ = _0051_ & _1112_;
  assign _0894_ = _0047_ & _1112_;
  assign _0896_ = _0061_ & _1112_;
  assign _0898_ = _0049_ & _1112_;
  assign _0649_ = _0053_ & _1116_;
  assign _0909_ = _0041_ & _1206_;
  assign _0912_ = 2'h0 & _1209_;
  assign _0916_ = 3'h0 & _1212_;
  assign _0960_ = _0485_ | _0486_;
  assign _0963_ = _0488_ | _0489_;
  assign _0966_ = _0491_ | _0492_;
  assign _0969_ = _0494_ | _0495_;
  assign _0972_ = _0497_ | _0498_;
  assign _0975_ = _0500_ | _0501_;
  assign _0978_ = _0503_ | _0504_;
  assign _0981_ = _0506_ | _0507_;
  assign _0984_ = _0509_ | _0510_;
  assign _0987_ = _0512_ | _0513_;
  assign _0990_ = _0515_ | _0516_;
  assign _0993_ = _0518_ | _0519_;
  assign _0999_ = _0524_ | _0525_;
  assign _1002_ = _0527_ | _0528_;
  assign _1005_ = _0530_ | _0531_;
  assign _1008_ = _0533_ | _0534_;
  assign _1009_ = _0536_ | _0516_;
  assign _0996_ = _0521_ | _0522_;
  assign _1015_ = _0542_ | _0543_;
  assign _1018_ = _0545_ | _0546_;
  assign _1024_ = _0552_ | _0553_;
  assign _1027_ = _0555_ | _0556_;
  assign _1030_ = _0558_ | _0559_;
  assign _1033_ = _0561_ | _0562_;
  assign _1036_ = _0564_ | _0565_;
  assign _1039_ = _0567_ | _0568_;
  assign _1042_ = _0570_ | _0571_;
  assign _1045_ = _0573_ | _0574_;
  assign _1048_ = _0576_ | _0577_;
  assign _1051_ = _0579_ | _0580_;
  assign _1054_ = _0582_ | _0583_;
  assign _1057_ = _0585_ | _0586_;
  assign _1060_ = _0588_ | _0589_;
  assign _1063_ = _0591_ | _0592_;
  assign _1066_ = _0594_ | _0595_;
  assign _1069_ = _0597_ | _0598_;
  assign _1072_ = _0600_ | _0601_;
  assign _1075_ = _0603_ | _0604_;
  assign _1078_ = _0606_ | _0607_;
  assign _1081_ = _0609_ | _0610_;
  assign _1084_ = _0612_ | _0613_;
  assign _1087_ = _0615_ | _0616_;
  assign _1090_ = _0618_ | _0619_;
  assign _1093_ = _0621_ | _0622_;
  assign _1096_ = _0624_ | _0625_;
  assign _1099_ = _0627_ | _0628_;
  assign _1103_ = _0632_ | _0633_;
  assign _1106_ = _0635_ | _0636_;
  assign _1109_ = _0638_ | _0639_;
  assign _1110_ = _0641_ | _0610_;
  assign _1113_ = _0643_ | _0644_;
  assign _1117_ = _0648_ | _0649_;
  assign _1118_ = _0651_ | _0652_;
  assign _1119_ = _0654_ | _0655_;
  assign _1123_ = _0659_ | _0660_;
  assign _1126_ = _0662_ | _0663_;
  assign _1129_ = _0665_ | _0666_;
  assign _1133_ = _0670_ | _0671_;
  assign _1136_ = _0673_ | _0674_;
  assign _1139_ = _0676_ | _0677_;
  assign _1140_ = _0679_ | _0680_;
  assign _1146_ = _0701_ | _0702_;
  assign _1149_ = _0704_ | _0705_;
  assign _1150_ = _0707_ | _0705_;
  assign _1012_ = _0539_ | _0540_;
  assign _1153_ = _0710_ | _0711_;
  assign _1157_ = _0734_ | _0735_;
  assign _1160_ = _0737_ | _0738_;
  assign _1163_ = _0740_ | _0741_;
  assign _1166_ = _0746_ | _0747_;
  assign _1169_ = _0749_ | _0750_;
  assign _1172_ = _0752_ | _0753_;
  assign _1175_ = _0755_ | _0756_;
  assign _1178_ = _0769_ | _0770_;
  assign _1185_ = _0809_ | _0810_;
  assign _1188_ = _0824_ | _0825_;
  assign _1192_ = _0849_ | _0850_;
  assign _1193_ = _0852_ | _0850_;
  assign _1200_ = _0881_ | _0882_;
  assign _1203_ = _0884_ | _0885_;
  assign _1204_ = _0884_ | _0887_;
  assign _1207_ = _0908_ | _0909_;
  assign _1210_ = _0911_ | _0912_;
  assign _1213_ = _0915_ | _0916_;
  assign _1214_ = _1342_ ^ 6'h09;
  assign _1215_ = _1344_ ^ _1340_;
  assign _1216_ = _1350_ ^ 6'h25;
  assign _1217_ = _1352_ ^ _1348_;
  assign _1218_ = _1354_ ^ _1346_;
  assign _1219_ = 6'h0a ^ _0126_;
  assign _1220_ = _1358_ ^ _1356_;
  assign _1221_ = _1364_ ^ _1362_;
  assign _1222_ = _1366_ ^ _1360_;
  assign _1223_ = _1368_ ^ 6'h16;
  assign _1224_ = _1374_ ^ _1372_;
  assign _1225_ = _1376_ ^ _1370_;
  assign _1226_ = _1380_ ^ _1378_;
  assign _1227_ = _1382_ ^ _0118_;
  assign _1228_ = 2'h3 ^ _0097_;
  assign _1229_ = _1386_ ^ 2'h2;
  assign _1230_ = _1388_ ^ _1384_;
  assign _1231_ = _0120_ ^ _0002_;
  assign _1232_ = _1390_ ^ _0008_;
  assign _1233_ = 6'h26 ^ _0110_;
  assign _1235_ = _1395_ ^ _1392_;
  assign _1236_ = _0116_ ^ 3'h3;
  assign _1237_ = _1399_ ^ _0105_;
  assign _1238_ = _1401_ ^ _1397_;
  assign _1239_ = _0102_ ^ _0112_;
  assign _1240_ = _1405_ ^ _1403_;
  assign _1241_ = _1409_ ^ _1407_;
  assign _1242_ = _1411_ ^ 2'h3;
  assign _1243_ = _1415_ ^ _1413_;
  assign _1244_ = _1417_ ^ _0006_;
  assign _1245_ = _1419_ ^ _0104_;
  assign _1246_ = _1420_ ^ 2'h1;
  assign _1247_ = _1422_ ^ _0038_;
  assign _1248_ = _1423_ ^ _0052_;
  assign _1249_ = _1425_ ^ _0057_;
  assign _1250_ = _0030_ ^ _0032_;
  assign _1251_ = _1428_ ^ _0012_;
  assign _1252_ = _1430_ ^ _1426_;
  assign _1253_ = _0114_ ^ _0122_;
  assign _1254_ = _1436_ ^ _0084_;
  assign _1255_ = _1438_ ^ _1434_;
  assign _1256_ = _1440_ ^ _1432_;
  assign _1257_ = _1442_ ^ _0068_;
  assign _1258_ = _0004_ ^ 6'h26;
  assign _1259_ = _0000_ ^ 6'h09;
  assign _1260_ = _0072_ ^ _0036_;
  assign _0487_ = { _0156_, _0156_, _0156_, _0156_, _0156_, _0156_ } & 6'h08;
  assign _0490_ = { _1494_, _1494_, _1494_, _1494_, _1494_, _1494_ } & 6'h0e;
  assign _0493_ = { _1492_, _1492_, _1492_, _1492_, _1492_, _1492_ } & _1214_;
  assign _0496_ = { _0923_, _0923_, _0923_, _0923_, _0923_, _0923_ } & _1215_;
  assign _0499_ = { _1498_, _1498_, _1498_, _1498_, _1498_, _1498_ } & 6'h01;
  assign _0502_ = { _1504_, _1504_, _1504_, _1504_, _1504_, _1504_ } & 6'h27;
  assign _0505_ = { _1502_, _1502_, _1502_, _1502_, _1502_, _1502_ } & _1216_;
  assign _0508_ = { _0925_, _0925_, _0925_, _0925_, _0925_, _0925_ } & _1217_;
  assign _0511_ = { _0324_, _0324_, _0324_, _0324_, _0324_, _0324_ } & _1218_;
  assign _0514_ = { _1510_, _1510_, _1510_, _1510_, _1510_, _1510_ } & _1219_;
  assign _0517_ = { _1514_, _1514_, _1514_, _1514_, _1514_, _1514_ } & 6'h07;
  assign _0520_ = { _0927_, _0927_, _0927_, _0927_, _0927_, _0927_ } & _1220_;
  assign _0523_ = { _1518_, _1518_, _1518_, _1518_, _1518_, _1518_ } & 6'h24;
  assign _0526_ = { _1522_, _1522_, _1522_, _1522_, _1522_, _1522_ } & 6'h25;
  assign _0529_ = { _0929_, _0929_, _0929_, _0929_, _0929_, _0929_ } & _1221_;
  assign _0532_ = { _0326_, _0326_, _0326_, _0326_, _0326_, _0326_ } & _1222_;
  assign _0535_ = { _1516_, _1516_, _1516_, _1516_, _1516_, _1516_ } & 6'h01;
  assign _0537_ = { _1514_, _1514_, _1514_, _1514_, _1514_, _1514_ } & _1223_;
  assign _0538_ = { _1518_, _1518_, _1518_, _1518_, _1518_, _1518_ } & 6'h0b;
  assign _0541_ = { _0056_, _0056_, _0056_, _0056_, _0056_, _0056_ } & 6'h31;
  assign _0544_ = { _0931_, _0931_, _0931_, _0931_, _0931_, _0931_ } & _1224_;
  assign _0547_ = { _0328_, _0328_, _0328_, _0328_, _0328_, _0328_ } & _1225_;
  assign _0549_ = _1508_ & _0109_;
  assign _0551_ = _1526_ & instr_first_cycle_i;
  assign _0554_ = _0933_ & _1226_;
  assign _0557_ = { _1472_, _1472_ } & _0107_;
  assign _0560_ = { _1468_, _1468_ } & _1227_;
  assign _0563_ = { _1526_, _1526_ } & _1228_;
  assign _0566_ = { _0136_, _0136_ } & _1229_;
  assign _0569_ = { _0330_, _0330_ } & _1230_;
  assign _0572_ = { _1508_, _1508_, _1508_, _1508_, _1508_, _1508_ } & _1231_;
  assign _0575_ = { _1472_, _1472_, _1472_, _1472_, _1472_, _1472_ } & _1232_;
  assign _0578_ = { _1526_, _1526_, _1526_, _1526_, _1526_, _1526_ } & _1233_;
  assign _0581_ = { _0167_, _0167_, _0167_, _0167_, _0167_, _0167_ } & _1234_;
  assign _0584_ = { _0332_, _0332_, _0332_, _0332_, _0332_, _0332_ } & _1235_;
  assign _0587_ = { _0158_, _0158_, _0158_ } & _1236_;
  assign _0590_ = { _0160_, _0160_, _0160_ } & 3'h5;
  assign _0593_ = { _1526_, _1526_, _1526_ } & _1237_;
  assign _0596_ = { _0935_, _0935_, _0935_ } & _1238_;
  assign _0599_ = { _1472_, _1472_, _1472_ } & _1239_;
  assign _0602_ = { _1530_, _1530_, _1530_ } & 3'h4;
  assign _0605_ = { _0937_, _0937_, _0937_ } & _1240_;
  assign _0608_ = { _1538_, _1538_ } & 2'h1;
  assign _0611_ = { _1542_, _1542_ } & 2'h1;
  assign _0614_ = { _0939_, _0939_ } & _1241_;
  assign _0617_ = { _1564_, _1564_ } & 2'h1;
  assign _0620_ = { _0153_, _0153_ } & _1242_;
  assign _0623_ = { _0144_, _0144_ } & 2'h1;
  assign _0626_ = { _0148_, _0148_ } & 2'h1;
  assign _0629_ = { _0941_, _0941_ } & _1243_;
  assign _0631_ = _0058_ & _0130_;
  assign _0634_ = _1574_ & _1244_;
  assign _0637_ = _1540_ & _1245_;
  assign _0640_ = { _1586_, _1586_ } & 2'h2;
  assign _0642_ = { _1542_, _1542_ } & _1246_;
  assign _0645_ = _1544_ & _1247_;
  assign _0647_ = _0133_ & _0059_;
  assign _0650_ = _1552_ & _1248_;
  assign _0653_ = _1552_ & _1249_;
  assign _0656_ = _1544_ & _1250_;
  assign _0658_ = _1576_ & _0128_;
  assign _0661_ = _1572_ & _1251_;
  assign _0664_ = _0943_ & _1252_;
  assign _0667_ = _1584_ & _1253_;
  assign _0669_ = _1591_ & _0320_;
  assign _0672_ = _0015_ & _1254_;
  assign _0675_ = _0945_ & _1255_;
  assign _0678_ = _0334_ & _1256_;
  assign _0681_ = _1544_ & _1257_;
  assign _0703_ = { instr_rdata_alu_i_t0[14], instr_rdata_alu_i_t0[14] } & 2'h3;
  assign _0706_ = { _0056_, _0056_ } & _0124_;
  assign _0708_ = { _0056_, _0056_ } & 2'h3;
  assign _0709_ = { _0056_, _0056_, _0056_, _0056_, _0056_, _0056_ } & 6'h26;
  assign _0712_ = { _1470_, _1470_, _1470_ } & 3'h5;
  assign _0731_ = instr_rdata_alu_i_t0[26] & _0076_;
  assign _0733_ = instr_rdata_alu_i_t0[26] & _0088_;
  assign _0736_ = { instr_rdata_alu_i_t0[26], instr_rdata_alu_i_t0[26], instr_rdata_alu_i_t0[26], instr_rdata_alu_i_t0[26], instr_rdata_alu_i_t0[26], instr_rdata_alu_i_t0[26] } & _1258_;
  assign _0739_ = { _1455_, _1455_, _1455_, _1455_, _1455_, _1455_ } & 6'h2e;
  assign _0742_ = { _1453_, _1453_, _1453_, _1453_, _1453_, _1453_ } & _1259_;
  assign _0748_ = { instr_rdata_alu_i_t0[14], instr_rdata_alu_i_t0[14], instr_rdata_alu_i_t0[14] } & 3'h1;
  assign _0751_ = { instr_first_cycle_i_t0, instr_first_cycle_i_t0 } & 2'h2;
  assign _0754_ = { instr_first_cycle_i_t0, instr_first_cycle_i_t0, instr_first_cycle_i_t0, instr_first_cycle_i_t0, instr_first_cycle_i_t0, instr_first_cycle_i_t0 } & _0100_;
  assign _0757_ = { instr_first_cycle_i_t0, instr_first_cycle_i_t0, instr_first_cycle_i_t0 } & _0102_;
  assign _0771_ = { _1528_, _1528_ } & 2'h2;
  assign _0777_ = _1508_ & _0044_;
  assign _0779_ = _1508_ & _0062_;
  assign _0782_ = _1468_ & _0321_;
  assign _0785_ = illegal_insn_o_t0 & rf_wdata_sel_o;
  assign _0787_ = illegal_insn_o_t0 & _0014_;
  assign _0789_ = illegal_insn_o_t0 & _0024_;
  assign _0791_ = illegal_insn_o_t0 & _0022_;
  assign _0793_ = illegal_insn_o_t0 & _0018_;
  assign _0795_ = illegal_insn_o_t0 & _0016_;
  assign _0797_ = illegal_insn_o_t0 & _0026_;
  assign _0799_ = illegal_c_insn_i_t0 & _0322_;
  assign _0803_ = _1462_ & _0139_;
  assign _0811_ = _0039_ & _1260_;
  assign _0813_ = _0039_ & _0095_;
  assign _0815_ = _0039_ & _0082_;
  assign _0817_ = _0039_ & _0078_;
  assign _0819_ = _0039_ & _0086_;
  assign _0821_ = _0039_ & _0080_;
  assign _0823_ = _0039_ & _0094_;
  assign _0826_ = { _0039_, _0039_ } & _0074_;
  assign _0828_ = _0058_ & _0059_;
  assign _0848_ = _1450_ & _0165_;
  assign _0851_ = { _1450_, _1450_ } & _0092_;
  assign _0853_ = { _1450_, _1450_ } & _0090_;
  assign _0855_ = _1580_ & _0318_;
  assign _0860_ = instr_rdata_i_t0[26] & _0319_;
  assign _0863_ = _1578_[0] & _0318_;
  assign _0865_ = _0150_ & _0317_;
  assign _0880_ = _1584_ & _0298_;
  assign _0883_ = { _0017_, _0017_ } & _0042_;
  assign _0886_ = { _1572_, _1572_ } & _0066_;
  assign _0888_ = { _1572_, _1572_ } & _0064_;
  assign _0889_ = _1544_ & _0038_;
  assign _0891_ = _1544_ & _0070_;
  assign _0893_ = _1544_ & _0050_;
  assign _0895_ = _1544_ & _0046_;
  assign _0897_ = _1544_ & _0060_;
  assign _0899_ = _1544_ & _0048_;
  assign _0907_ = _1552_ & _0052_;
  assign _0910_ = { _1544_, _1544_ } & _0040_;
  assign _0913_ = { _1458_, _1458_ } & csr_op;
  assign _0917_ = { branch_taken_i_t0, branch_taken_i_t0, branch_taken_i_t0 } & 3'h7;
  assign _0919_ = illegal_insn_o_t0 & mult_sel_o;
  assign _0921_ = illegal_insn_o_t0 & div_sel_o;
  assign _1341_ = _0487_ | _0960_;
  assign _1343_ = _0490_ | _0963_;
  assign _1345_ = _0493_ | _0966_;
  assign _1347_ = _0496_ | _0969_;
  assign _1349_ = _0499_ | _0972_;
  assign _1351_ = _0502_ | _0975_;
  assign _1353_ = _0505_ | _0978_;
  assign _1355_ = _0508_ | _0981_;
  assign _0005_ = _0511_ | _0984_;
  assign _1357_ = _0514_ | _0987_;
  assign _1359_ = _0517_ | _0990_;
  assign _1361_ = _0520_ | _0993_;
  assign _1363_ = _0523_ | _0996_;
  assign _1365_ = _0526_ | _0999_;
  assign _1367_ = _0529_ | _1002_;
  assign _0121_ = _0532_ | _1005_;
  assign _1369_ = _0535_ | _1008_;
  assign _1371_ = _0537_ | _1009_;
  assign _1373_ = _0538_ | _0996_;
  assign _1375_ = _0541_ | _1012_;
  assign _1377_ = _0544_ | _1015_;
  assign _0101_ = _0547_ | _1018_;
  assign _1379_ = _0549_ | _0548_;
  assign _1381_ = _0551_ | _0550_;
  assign alu_op_b_mux_sel_o_t0 = _0554_ | _1024_;
  assign _1383_ = _0557_ | _1027_;
  assign _1385_ = _0560_ | _1030_;
  assign _1387_ = _0563_ | _1033_;
  assign _1389_ = _0566_ | _1036_;
  assign alu_op_a_mux_sel_o_t0 = _0569_ | _1039_;
  assign _1391_ = _0572_ | _1042_;
  assign _1393_ = _0575_ | _1045_;
  assign _1394_ = _0578_ | _1048_;
  assign _1396_ = _0581_ | _1051_;
  assign alu_operator_o_t0 = _0584_ | _1054_;
  assign _1398_ = _0587_ | _1057_;
  assign _1400_ = _0590_ | _1060_;
  assign _1402_ = _0593_ | _1063_;
  assign imm_b_mux_sel_o_t0 = _0596_ | _1066_;
  assign _1404_ = _0599_ | _1069_;
  assign _1406_ = _0602_ | _1072_;
  assign bt_b_mux_sel_o_t0 = _0605_ | _1075_;
  assign _1408_ = _0608_ | _1078_;
  assign _1410_ = _0611_ | _1081_;
  assign _0075_ = _0614_ | _1084_;
  assign _1412_ = _0617_ | _1087_;
  assign _0093_ = _0620_ | _1090_;
  assign _1414_ = _0623_ | _1093_;
  assign _1416_ = _0626_ | _1096_;
  assign _0091_ = _0629_ | _1099_;
  assign _1418_ = _0631_ | _0630_;
  assign _0129_ = _0634_ | _1103_;
  assign _0123_ = _0637_ | _1106_;
  assign _1421_ = _0640_ | _1109_;
  assign _0043_ = _0642_ | _1110_;
  assign _0027_ = _0645_ | _1113_;
  assign _1424_ = _0647_ | _0646_;
  assign _0025_ = _0650_ | _1117_;
  assign _0023_ = _0653_ | _1118_;
  assign _1427_ = _0656_ | _1119_;
  assign _1429_ = _0658_ | _0657_;
  assign _1431_ = _0661_ | _1123_;
  assign _1433_ = _0664_ | _1126_;
  assign _1435_ = _0667_ | _1129_;
  assign _1437_ = _0669_ | _0668_;
  assign _1439_ = _0672_ | _1133_;
  assign _1441_ = _0675_ | _1136_;
  assign _0021_ = _0678_ | _1139_;
  assign rf_ren_a_o_t0 = _0681_ | _1140_;
  assign _0125_ = _0703_ | _1146_;
  assign _0119_ = _0706_ | _1149_;
  assign _0108_ = _0708_ | _1150_;
  assign _0009_ = _0709_ | _1012_;
  assign _0113_ = _0712_ | _1153_;
  assign _0045_ = _0731_ | _0730_;
  assign _0063_ = _0733_ | _0732_;
  assign _0003_ = _0736_ | _1157_;
  assign _0001_ = _0739_ | _1160_;
  assign _0127_ = _0742_ | _1163_;
  assign _0117_ = _0748_ | _1166_;
  assign _0098_ = _0751_ | _1169_;
  assign _0111_ = _0754_ | _1172_;
  assign _0106_ = _0757_ | _1175_;
  assign bt_a_mux_sel_o_t0 = _0771_ | _1178_;
  assign div_sel_o_t0 = _0777_ | _0776_;
  assign mult_sel_o_t0 = _0779_ | _0778_;
  assign imm_a_mux_sel_o_t0 = _0782_ | _0781_;
  assign csr_access_o_t0 = _0785_ | _0784_;
  assign branch_in_dec_o_t0 = _0787_ | _0786_;
  assign jump_set_o_t0 = _0789_ | _0788_;
  assign jump_in_dec_o_t0 = _0791_ | _0790_;
  assign data_we_o_t0 = _0793_ | _0792_;
  assign data_req_o_t0 = _0795_ | _0794_;
  assign rf_we_o_t0 = _0797_ | _0796_;
  assign illegal_insn_o_t0 = _0799_ | _0798_;
  assign _0037_ = _0803_ | _0802_;
  assign _0033_ = _0811_ | _1185_;
  assign _0071_ = _0813_ | _0812_;
  assign _0051_ = _0815_ | _0814_;
  assign _0047_ = _0817_ | _0816_;
  assign _0061_ = _0819_ | _0818_;
  assign _0049_ = _0821_ | _0820_;
  assign _0069_ = _0823_ | _0822_;
  assign _0041_ = _0826_ | _1188_;
  assign _0053_ = _0828_ | _0827_;
  assign _0013_ = _0848_ | _0847_;
  assign _0067_ = _0851_ | _1192_;
  assign _0065_ = _0853_ | _1193_;
  assign _0011_ = _0855_ | _0854_;
  assign _0007_ = _0860_ | _0859_;
  assign _0131_ = _0863_ | _0862_;
  assign _0115_ = _0865_ | _0864_;
  assign data_sign_extension_o_t0 = _0880_ | _0879_;
  assign data_type_o_t0 = _0883_ | _1200_;
  assign multdiv_signed_mode_o_t0 = _0886_ | _1203_;
  assign multdiv_operator_o_t0 = _0888_ | _1204_;
  assign rf_wdata_sel_o_t0 = _0889_ | _0644_;
  assign wfi_insn_o_t0 = _0891_ | _0890_;
  assign ecall_insn_o_t0 = _0893_ | _0892_;
  assign dret_insn_o_t0 = _0895_ | _0894_;
  assign mret_insn_o_t0 = _0897_ | _0896_;
  assign ebrk_insn_o_t0 = _0899_ | _0898_;
  assign icache_inval_o_t0 = _0907_ | _0649_;
  assign csr_op_t0 = _0910_ | _1207_;
  assign csr_op_o_t0 = _0913_ | _1210_;
  assign _0103_ = _0917_ | _1213_;
  assign mult_en_o_t0 = _0919_ | _0918_;
  assign div_en_o_t0 = _0921_ | _0920_;
  assign _0317_ = ~ _0104_;
  assign _0319_ = ~ _0010_;
  assign _0320_ = ~ _0054_;
  assign _0321_ = ~ _0055_;
  assign _0322_ = ~ _0020_;
  assign _0132_ = | { _1592_, _1590_ };
  assign _0134_ = | { _1587_, _1583_ };
  assign _0135_ = | { _1531_, _1529_, _1527_ };
  assign _0137_ = | { _1550_, _1451_ };
  assign _0138_ = | { _1589_, _1587_, _1571_ };
  assign _0139_ = | { _1549_, _1548_, _1547_, _1546_, _1545_ };
  assign _0141_ = | { _1596_, _1594_, _1592_, _1590_, _1575_, _1571_ };
  assign _0143_ = | { _1555_, _1553_ };
  assign _0145_ = | { _1559_, _1557_ };
  assign _0147_ = | { _1565_, _1563_, _1561_ };
  assign _0151_ = | { _1487_, _1485_, _1483_, _1481_ };
  assign _0152_ = | { _1565_, _1559_, _1555_ };
  assign _0154_ = | { _1479_, _1477_, _1475_, _1473_ };
  assign _0155_ = | { _1505_, _1487_, _1485_, _1483_, _1481_, _1479_, _1477_, _1475_, _1473_ };
  assign _0157_ = | { _1535_, _1531_ };
  assign _0159_ = | { _1529_, _1527_ };
  assign _0161_ = | { _1590_, _1589_, _1587_, _1583_, _1575_, _1571_ };
  assign _0165_ = | { _1569_, _1567_, _1565_, _1563_, _1561_, _1559_, _1557_, _1555_, _1553_ };
  assign _0166_ = | { _1535_, _1533_, _1531_, _1529_, _1527_, _1523_ };
  assign _0190_ = ~ _1489_;
  assign _0192_ = ~ _1499_;
  assign _0196_ = ~ _1519_;
  assign _0194_ = ~ _1469_;
  assign _0198_ = ~ _1523_;
  assign _0205_ = ~ _0145_;
  assign _0191_ = ~ _0155_;
  assign _0193_ = ~ _1497_;
  assign _0195_ = ~ _1509_;
  assign _0197_ = ~ _1517_;
  assign _0200_ = ~ _0157_;
  assign _0202_ = ~ _1471_;
  assign _0204_ = ~ _1537_;
  assign _0206_ = ~ _0143_;
  assign _0443_ = _1490_ & _0191_;
  assign _0446_ = _1500_ & _0193_;
  assign _0449_ = _1470_ & _0195_;
  assign _0452_ = _1520_ & _0197_;
  assign _0455_ = _1470_ & _0197_;
  assign _0458_ = _1524_ & _0199_;
  assign _0461_ = _1524_ & _0200_;
  assign _0464_ = _1526_ & _0202_;
  assign _0467_ = _1540_ & _0204_;
  assign _0470_ = _0146_ & _0206_;
  assign _0473_ = _1552_ & _0208_;
  assign _0476_ = _0019_ & _0210_;
  assign _0444_ = _0156_ & _0190_;
  assign _0447_ = _1498_ & _0192_;
  assign _0450_ = _1510_ & _0194_;
  assign _0453_ = _1518_ & _0196_;
  assign _0456_ = _1518_ & _0194_;
  assign _0459_ = _1508_ & _0198_;
  assign _0462_ = _0158_ & _0198_;
  assign _0465_ = _1472_ & _0201_;
  assign _0468_ = _1538_ & _0203_;
  assign _0471_ = _0144_ & _0205_;
  assign _0474_ = _1544_ & _0207_;
  assign _0477_ = _1584_ & _0209_;
  assign _0445_ = _1490_ & _0156_;
  assign _0448_ = _1500_ & _1498_;
  assign _0451_ = _1470_ & _1510_;
  assign _0454_ = _1520_ & _1518_;
  assign _0457_ = _1470_ & _1518_;
  assign _0460_ = _1524_ & _1508_;
  assign _0463_ = _1524_ & _0158_;
  assign _0466_ = _1526_ & _1472_;
  assign _0469_ = _1540_ & _1538_;
  assign _0472_ = _0146_ & _0144_;
  assign _0475_ = _1552_ & _1544_;
  assign _0478_ = _0019_ & _1584_;
  assign _0946_ = _0443_ | _0444_;
  assign _0947_ = _0446_ | _0447_;
  assign _0948_ = _0449_ | _0450_;
  assign _0949_ = _0452_ | _0453_;
  assign _0950_ = _0455_ | _0456_;
  assign _0951_ = _0458_ | _0459_;
  assign _0952_ = _0461_ | _0462_;
  assign _0953_ = _0464_ | _0465_;
  assign _0954_ = _0467_ | _0468_;
  assign _0955_ = _0470_ | _0471_;
  assign _0956_ = _0473_ | _0474_;
  assign _0957_ = _0476_ | _0477_;
  assign _0923_ = _0946_ | _0445_;
  assign _0925_ = _0947_ | _0448_;
  assign _0927_ = _0948_ | _0451_;
  assign _0929_ = _0949_ | _0454_;
  assign _0931_ = _0950_ | _0457_;
  assign _0933_ = _0951_ | _0460_;
  assign _0935_ = _0952_ | _0463_;
  assign _0937_ = _0953_ | _0466_;
  assign _0939_ = _0954_ | _0469_;
  assign _0941_ = _0955_ | _0472_;
  assign _0943_ = _0956_ | _0475_;
  assign _0945_ = _0957_ | _0478_;
  assign _0140_ = | { _1541_, _1539_, _1537_ };
  assign _0149_ = | { _1585_, _1541_, _1539_ };
  assign _0163_ = | { _1585_, _1541_ };
  assign _0922_ = _1489_ | _0155_;
  assign _0924_ = _1499_ | _1497_;
  assign _0926_ = _1469_ | _1509_;
  assign _0928_ = _1519_ | _1517_;
  assign _0930_ = _1469_ | _1517_;
  assign _0932_ = _1523_ | _1507_;
  assign _0934_ = _1523_ | _0157_;
  assign _0936_ = _1525_ | _1471_;
  assign _0938_ = _1539_ | _1537_;
  assign _0940_ = _0145_ | _0143_;
  assign _0942_ = _1551_ | _1543_;
  assign _0944_ = _1587_ | _1583_;
  assign _0323_ = | { _0922_, _1495_, _1493_, _1491_ };
  assign _0325_ = | { _1515_, _1513_, _0926_ };
  assign _0327_ = | { _1515_, _1513_, _1509_ };
  assign _0329_ = | { _1533_, _1523_, _1511_, _1507_, _1471_, _1467_ };
  assign _0331_ = | { _1511_, _1507_, _1471_ };
  assign _0333_ = | { _0942_, _1596_, _1594_, _1592_, _1575_, _1571_ };
  assign _1340_ = _0155_ ? 6'h00 : 6'h08;
  assign _1342_ = _1493_ ? 6'h0a : 6'h04;
  assign _1344_ = _1491_ ? 6'h09 : _1342_;
  assign _1346_ = _0922_ ? _1340_ : _1344_;
  assign _1348_ = _1497_ ? 6'h03 : 6'h02;
  assign _1350_ = _1503_ ? 6'h01 : 6'h26;
  assign _1352_ = _1501_ ? 6'h25 : _1350_;
  assign _1354_ = _0924_ ? _1348_ : _1352_;
  assign _0004_ = _0323_ ? _1346_ : _1354_;
  assign _1356_ = _1509_ ? _0126_ : 6'h0a;
  assign _1358_ = _1513_ ? 6'h04 : 6'h03;
  assign _1360_ = _0926_ ? _1356_ : _1358_;
  assign _1362_ = _1517_ ? 6'h02 : 6'h26;
  assign _1364_ = _1521_ ? 6'h25 : 6'h00;
  assign _1366_ = _0928_ ? _1362_ : _1364_;
  assign _0120_ = _0325_ ? _1360_ : _1366_;
  assign _1368_ = _1515_ ? 6'h14 : 6'h15;
  assign _1370_ = _1513_ ? 6'h16 : _1368_;
  assign _1372_ = _1517_ ? 6'h13 : 6'h18;
  assign _1374_ = _1456_ ? 6'h17 : 6'h26;
  assign _1376_ = _0930_ ? _1372_ : _1374_;
  assign _0100_ = _0327_ ? _1370_ : _1376_;
  assign _1378_ = _1507_ ? 1'h0 : _0109_;
  assign _1380_ = _1525_ ? _0099_ : 1'h1;
  assign alu_op_b_mux_sel_o = _0932_ ? _1378_ : _1380_;
  assign _1382_ = _1471_ ? _0107_ : 2'h0;
  assign _1384_ = _1467_ ? _0118_ : _1382_;
  assign _1386_ = _1525_ ? _0097_ : 2'h3;
  assign _1388_ = _0135_ ? 2'h2 : _1386_;
  assign alu_op_a_mux_sel_o = _0329_ ? _1384_ : _1388_;
  assign _1390_ = _1507_ ? _0002_ : _0120_;
  assign _1392_ = _1471_ ? _0008_ : _1390_;
  assign _1234_ = _1525_ ? _0110_ : 6'h26;
  assign _1395_ = _0166_ ? 6'h00 : _1234_;
  assign alu_operator_o = _0331_ ? _1392_ : _1395_;
  assign _1397_ = _0157_ ? 3'h3 : _0116_;
  assign _1399_ = _0159_ ? 3'h5 : 3'h0;
  assign _1401_ = _1525_ ? _0105_ : _1399_;
  assign imm_b_mux_sel_o = _0934_ ? _1397_ : _1401_;
  assign _1403_ = _1471_ ? _0112_ : _0102_;
  assign _1405_ = _1529_ ? 3'h4 : 3'h0;
  assign bt_b_mux_sel_o = _0936_ ? _1403_ : _1405_;
  assign _1407_ = _1537_ ? 2'h3 : 2'h2;
  assign _1409_ = _1541_ ? 2'h1 : 2'h0;
  assign _0074_ = _0938_ ? _1407_ : _1409_;
  assign _1411_ = _1563_ ? 2'h1 : 2'h0;
  assign _0092_ = _0152_ ? 2'h3 : _1411_;
  assign _1413_ = _0143_ ? 2'h3 : 2'h2;
  assign _1415_ = _0147_ ? 2'h1 : 2'h0;
  assign _0090_ = _0940_ ? _1413_ : _1415_;
  assign _1417_ = _1550_ ? _0130_ : 1'h0;
  assign _0128_ = _1573_ ? _0006_ : _1417_;
  assign _1419_ = _0163_ ? 1'h0 : 1'h1;
  assign _0122_ = _1539_ ? _0104_ : _1419_;
  assign _1420_ = _1585_ ? 2'h2 : 2'h0;
  assign _0042_ = _1541_ ? 2'h1 : _1420_;
  assign _1422_ = _0141_ ? 1'h1 : 1'h0;
  assign _0026_ = _1543_ ? _0038_ : _1422_;
  assign _1423_ = _0132_ ? _0059_ : 1'h0;
  assign _0024_ = _1551_ ? _0052_ : _1423_;
  assign _1425_ = _0132_ ? 1'h1 : 1'h0;
  assign _0022_ = _1551_ ? _0057_ : _1425_;
  assign _1426_ = _1543_ ? _0032_ : _0030_;
  assign _1428_ = _1575_ ? _0128_ : 1'h0;
  assign _1430_ = _1571_ ? _0012_ : _1428_;
  assign _1432_ = _0942_ ? _1426_ : _1430_;
  assign _1434_ = _1583_ ? _0122_ : _0114_;
  assign _1436_ = _1590_ ? _0054_ : 1'h1;
  assign _1438_ = _1589_ ? _0084_ : _1436_;
  assign _1440_ = _0944_ ? _1434_ : _1438_;
  assign _0020_ = _0333_ ? _1432_ : _1440_;
  assign _1442_ = _0161_ ? 1'h1 : 1'h0;
  assign rf_ren_a_o = _1543_ ? _0068_ : _1442_;
  assign _1443_ = csr_op == 2'h2;
  assign _1445_ = csr_op == 2'h3;
  assign _1447_ = ! instr_rdata_i[19:15];
  assign _1449_ = { instr_rdata_i[26], instr_rdata_i[13:12] } == 3'h5;
  assign _1452_ = ! instr_rdata_alu_i[31:27];
  assign _1454_ = instr_rdata_alu_i[31:27] == 5'h08;
  assign _1457_ = _1459_ && _1447_;
  assign _1459_ = _1443_ || _1445_;
  assign _1461_ = _1464_ || _1465_;
  assign _1463_ = | instr_rdata_i[14:12];
  assign _1464_ = | instr_rdata_i[19:15];
  assign _1465_ = | instr_rdata_i[11:7];
  assign _0124_ = instr_rdata_alu_i[14] ? 2'h3 : 2'h0;
  assign _0118_ = _1456_ ? 2'h0 : _0124_;
  assign _0055_ = _1456_ ? 1'h1 : 1'h0;
  assign _0107_ = _1456_ ? 2'h0 : 2'h3;
  assign _0008_ = _1456_ ? 6'h00 : 6'h26;
  assign _0112_ = _1469_ ? 3'h5 : 3'h0;
  assign _1489_ = { instr_rdata_alu_i[31:25], instr_rdata_alu_i[14:12] } == 10'h105;
  assign _1491_ = { instr_rdata_alu_i[31:25], instr_rdata_alu_i[14:12] } == 10'h005;
  assign _1493_ = { instr_rdata_alu_i[31:25], instr_rdata_alu_i[14:12] } == 10'h001;
  assign _1495_ = { instr_rdata_alu_i[31:25], instr_rdata_alu_i[14:12] } == 10'h007;
  assign _1497_ = { instr_rdata_alu_i[31:25], instr_rdata_alu_i[14:12] } == 10'h006;
  assign _1499_ = { instr_rdata_alu_i[31:25], instr_rdata_alu_i[14:12] } == 10'h004;
  assign _1501_ = { instr_rdata_alu_i[31:25], instr_rdata_alu_i[14:12] } == 10'h002;
  assign _1503_ = { instr_rdata_alu_i[31:25], instr_rdata_alu_i[14:12] } == 10'h100;
  assign _1505_ = ! { instr_rdata_alu_i[31:25], instr_rdata_alu_i[14:12] };
  assign _0076_ = _0154_ ? 1'h1 : 1'h0;
  assign _1473_ = { instr_rdata_alu_i[31:25], instr_rdata_alu_i[14:12] } == 10'h00f;
  assign _1475_ = { instr_rdata_alu_i[31:25], instr_rdata_alu_i[14:12] } == 10'h00e;
  assign _1477_ = { instr_rdata_alu_i[31:25], instr_rdata_alu_i[14:12] } == 10'h00d;
  assign _1479_ = { instr_rdata_alu_i[31:25], instr_rdata_alu_i[14:12] } == 10'h00c;
  assign _0088_ = _0151_ ? 1'h1 : 1'h0;
  assign _1481_ = { instr_rdata_alu_i[31:25], instr_rdata_alu_i[14:12] } == 10'h00b;
  assign _1483_ = { instr_rdata_alu_i[31:25], instr_rdata_alu_i[14:12] } == 10'h00a;
  assign _1485_ = { instr_rdata_alu_i[31:25], instr_rdata_alu_i[14:12] } == 10'h009;
  assign _1487_ = { instr_rdata_alu_i[31:25], instr_rdata_alu_i[14:12] } == 10'h008;
  assign _0044_ = instr_rdata_alu_i[26] ? 1'h0 : _0076_;
  assign _0062_ = instr_rdata_alu_i[26] ? 1'h0 : _0088_;
  assign _0002_ = instr_rdata_alu_i[26] ? 6'h26 : _0004_;
  assign _0000_ = _1454_ ? 6'h08 : 6'h26;
  assign _0126_ = _1452_ ? 6'h09 : _0000_;
  assign _1519_ = instr_rdata_alu_i[14:12] == 3'h3;
  assign _1521_ = instr_rdata_alu_i[14:12] == 3'h2;
  assign _0109_ = instr_rdata_alu_i[14] ? 1'h0 : 1'h1;
  assign _0116_ = instr_rdata_alu_i[14] ? 3'h0 : 3'h1;
  assign _0099_ = instr_first_cycle_i ? 1'h0 : 1'h1;
  assign _0097_ = instr_first_cycle_i ? 2'h0 : 2'h2;
  assign _0110_ = instr_first_cycle_i ? _0100_ : 6'h00;
  assign _0105_ = instr_first_cycle_i ? 3'h0 : _0102_;
  assign _1513_ = instr_rdata_alu_i[14:12] == 3'h7;
  assign _1515_ = instr_rdata_alu_i[14:12] == 3'h6;
  assign _1509_ = instr_rdata_alu_i[14:12] == 3'h5;
  assign _1517_ = instr_rdata_alu_i[14:12] == 3'h4;
  assign _1469_ = instr_rdata_alu_i[14:12] == 3'h1;
  assign _1456_ = ! instr_rdata_alu_i[14:12];
  assign _1511_ = instr_rdata_alu_i[6:0] == 7'h13;
  assign _1533_ = instr_rdata_alu_i[6:0] == 7'h03;
  assign _1531_ = instr_rdata_alu_i[6:0] == 7'h17;
  assign _1535_ = instr_rdata_alu_i[6:0] == 7'h37;
  assign _1523_ = instr_rdata_alu_i[6:0] == 7'h23;
  assign bt_a_mux_sel_o = _1527_ ? 2'h0 : 2'h2;
  assign _1471_ = instr_rdata_alu_i[6:0] == 7'h0f;
  assign _1525_ = instr_rdata_alu_i[6:0] == 7'h63;
  assign _1527_ = instr_rdata_alu_i[6:0] == 7'h67;
  assign _1529_ = instr_rdata_alu_i[6:0] == 7'h6f;
  assign div_sel_o = _1507_ ? _0044_ : 1'h0;
  assign mult_sel_o = _1507_ ? _0062_ : 1'h0;
  assign _1507_ = instr_rdata_alu_i[6:0] == 7'h33;
  assign imm_a_mux_sel_o = _1467_ ? _0055_ : 1'h1;
  assign _1467_ = instr_rdata_alu_i[6:0] == 7'h73;
  assign csr_access_o = illegal_insn_o ? 1'h0 : rf_wdata_sel_o;
  assign branch_in_dec_o = illegal_insn_o ? 1'h0 : _0014_;
  assign jump_set_o = illegal_insn_o ? 1'h0 : _0024_;
  assign jump_in_dec_o = illegal_insn_o ? 1'h0 : _0022_;
  assign data_we_o = illegal_insn_o ? 1'h0 : _0018_;
  assign data_req_o = illegal_insn_o ? 1'h0 : _0016_;
  assign rf_we_o = illegal_insn_o ? 1'h0 : _0026_;
  assign illegal_insn_o = illegal_c_insn_i ? 1'h1 : _0020_;
  assign _0072_ = _0140_ ? 1'h0 : 1'h1;
  assign _1537_ = instr_rdata_i[13:12] == 2'h3;
  assign _0094_ = instr_rdata_i[14] ? 1'h0 : 1'h1;
  assign _0036_ = _1461_ ? 1'h1 : _0034_;
  assign _0082_ = _1545_ ? 1'h1 : 1'h0;
  assign _0034_ = _0139_ ? 1'h0 : 1'h1;
  assign _1545_ = ! instr_rdata_i[31:20];
  assign _0095_ = _1546_ ? 1'h1 : 1'h0;
  assign _1546_ = instr_rdata_i[31:20] == 12'h105;
  assign _0078_ = _1547_ ? 1'h1 : 1'h0;
  assign _1547_ = instr_rdata_i[31:20] == 12'h7b2;
  assign _0086_ = _1548_ ? 1'h1 : 1'h0;
  assign _1548_ = instr_rdata_i[31:20] == 12'h302;
  assign _0080_ = _1549_ ? 1'h1 : 1'h0;
  assign _1549_ = instr_rdata_i[31:20] == 12'h001;
  assign _0032_ = _1451_ ? _0036_ : _0072_;
  assign _0070_ = _1451_ ? _0095_ : 1'h0;
  assign _0050_ = _1451_ ? _0082_ : 1'h0;
  assign _0046_ = _1451_ ? _0078_ : 1'h0;
  assign _0060_ = _1451_ ? _0086_ : 1'h0;
  assign _0048_ = _1451_ ? _0080_ : 1'h0;
  assign _0038_ = _1451_ ? 1'h0 : 1'h1;
  assign _0068_ = _1451_ ? 1'h0 : _0094_;
  assign _0040_ = _1451_ ? 2'h0 : _0074_;
  assign _0059_ = instr_first_cycle_i ? 1'h1 : 1'h0;
  assign _0030_ = _0137_ ? 1'h0 : 1'h1;
  assign _0057_ = _1550_ ? 1'h1 : 1'h0;
  assign _0052_ = _1550_ ? _0059_ : 1'h0;
  assign _0028_ = _0165_ ? 1'h0 : 1'h1;
  assign _1567_ = { instr_rdata_i[31:25], instr_rdata_i[14:12] } == 10'h008;
  assign _1569_[0] = ! { instr_rdata_i[31:25], instr_rdata_i[14:12] };
  assign _1569_[1] = { instr_rdata_i[31:25], instr_rdata_i[14:12] } == 10'h100;
  assign _1569_[2] = { instr_rdata_i[31:25], instr_rdata_i[14:12] } == 10'h002;
  assign _1569_[3] = { instr_rdata_i[31:25], instr_rdata_i[14:12] } == 10'h003;
  assign _1569_[4] = { instr_rdata_i[31:25], instr_rdata_i[14:12] } == 10'h004;
  assign _1569_[5] = { instr_rdata_i[31:25], instr_rdata_i[14:12] } == 10'h006;
  assign _1569_[6] = { instr_rdata_i[31:25], instr_rdata_i[14:12] } == 10'h007;
  assign _1569_[7] = { instr_rdata_i[31:25], instr_rdata_i[14:12] } == 10'h001;
  assign _1569_[8] = { instr_rdata_i[31:25], instr_rdata_i[14:12] } == 10'h005;
  assign _1569_[9] = { instr_rdata_i[31:25], instr_rdata_i[14:12] } == 10'h105;
  assign _1553_ = { instr_rdata_i[31:25], instr_rdata_i[14:12] } == 10'h00f;
  assign _1555_ = { instr_rdata_i[31:25], instr_rdata_i[14:12] } == 10'h00e;
  assign _1557_ = { instr_rdata_i[31:25], instr_rdata_i[14:12] } == 10'h00d;
  assign _1559_ = { instr_rdata_i[31:25], instr_rdata_i[14:12] } == 10'h00c;
  assign _1561_ = { instr_rdata_i[31:25], instr_rdata_i[14:12] } == 10'h00b;
  assign _1563_ = { instr_rdata_i[31:25], instr_rdata_i[14:12] } == 10'h00a;
  assign _1565_ = { instr_rdata_i[31:25], instr_rdata_i[14:12] } == 10'h009;
  assign _0012_ = _1449_ ? 1'h1 : _0028_;
  assign _0066_ = _1449_ ? 2'h0 : _0092_;
  assign _0064_ = _1449_ ? 2'h0 : _0090_;
  assign _0010_ = _1579_ ? _1598_ : 1'h1;
  assign _1579_ = | _1577_;
  assign _1577_[1] = instr_rdata_i[31:27] == 5'h08;
  assign _0006_ = instr_rdata_i[26] ? 1'h1 : _0010_;
  assign _0318_ = ! instr_rdata_i[26:25];
  assign _0130_ = _1577_[0] ? _1598_ : 1'h1;
  assign _1577_[0] = ! instr_rdata_i[31:27];
  assign _0104_ = instr_rdata_i[14] ? 1'h1 : 1'h0;
  assign _0114_ = _0149_ ? _0104_ : 1'h1;
  assign _1539_ = instr_rdata_i[13:12] == 2'h2;
  assign _1541_ = instr_rdata_i[13:12] == 2'h1;
  assign _1585_ = ! instr_rdata_i[13:12];
  assign _0084_ = _1588_ ? 1'h0 : 1'h1;
  assign _1588_ = | { _1581_[5:3], _1573_, _1550_, _1451_ };
  assign _1451_ = ! instr_rdata_i[14:12];
  assign _1550_ = instr_rdata_i[14:12] == 3'h1;
  assign _1581_[3] = instr_rdata_i[14:12] == 3'h4;
  assign _1573_ = instr_rdata_i[14:12] == 3'h5;
  assign _1581_[4] = instr_rdata_i[14:12] == 3'h6;
  assign _1581_[5] = instr_rdata_i[14:12] == 3'h7;
  assign _0054_ = _1463_ ? 1'h1 : 1'h0;
  assign _1551_ = instr_rdata_i[6:0] == 7'h0f;
  assign _1594_ = instr_rdata_i[6:0] == 7'h17;
  assign _1596_ = instr_rdata_i[6:0] == 7'h37;
  assign _1592_ = instr_rdata_i[6:0] == 7'h6f;
  assign _0014_ = _1589_ ? 1'h1 : 1'h0;
  assign data_sign_extension_o = _1583_ ? _0298_ : 1'h0;
  assign data_type_o = _0134_ ? _0042_ : 2'h0;
  assign multdiv_signed_mode_o = _1571_ ? _0066_ : 2'h0;
  assign multdiv_operator_o = _1571_ ? _0064_ : 2'h0;
  assign rf_wdata_sel_o = _1543_ ? _0038_ : 1'h0;
  assign wfi_insn_o = _1543_ ? _0070_ : 1'h0;
  assign ecall_insn_o = _1543_ ? _0050_ : 1'h0;
  assign dret_insn_o = _1543_ ? _0046_ : 1'h0;
  assign mret_insn_o = _1543_ ? _0060_ : 1'h0;
  assign ebrk_insn_o = _1543_ ? _0048_ : 1'h0;
  assign rf_ren_b_o = _0138_ ? 1'h1 : 1'h0;
  assign _1571_ = instr_rdata_i[6:0] == 7'h33;
  assign _1575_ = instr_rdata_i[6:0] == 7'h13;
  assign _1583_ = instr_rdata_i[6:0] == 7'h03;
  assign _1587_ = instr_rdata_i[6:0] == 7'h23;
  assign _1589_ = instr_rdata_i[6:0] == 7'h63;
  assign _1590_ = instr_rdata_i[6:0] == 7'h67;
  assign _1543_ = instr_rdata_i[6:0] == 7'h73;
  assign icache_inval_o = _1551_ ? _0052_ : 1'h0;
  assign csr_op = _1543_ ? _0040_ : 2'h0;
  assign _0018_ = _1587_ ? 1'h1 : 1'h0;
  assign _0016_ = _0134_ ? 1'h1 : 1'h0;
  assign csr_op_o = _1457_ ? 2'h0 : csr_op;
  assign _1598_ = _0318_ ? 1'h0 : 1'h1;
  assign _0102_ = branch_taken_i ? 3'h2 : 3'h5;
  assign mult_en_o = illegal_insn_o ? 1'h0 : mult_sel_o;
  assign div_en_o = illegal_insn_o ? 1'h0 : div_sel_o;
  assign _1581_[0] = _1451_;
  assign _1582_[0] = _0039_;
  assign alu_multicycle_o = 1'h0;
  assign alu_multicycle_o_t0 = 1'h0;
  assign imm_b_type_o = { instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[7], instr_rdata_i[30:25], instr_rdata_i[11:8], 1'h0 };
  assign imm_b_type_o_t0 = { instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[7], instr_rdata_i_t0[30:25], instr_rdata_i_t0[11:8], 1'h0 };
  assign imm_i_type_o = { instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31:20] };
  assign imm_i_type_o_t0 = { instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31:20] };
  assign imm_j_type_o = { instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[19:12], instr_rdata_i[20], instr_rdata_i[30:21], 1'h0 };
  assign imm_j_type_o_t0 = { instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[19:12], instr_rdata_i_t0[20], instr_rdata_i_t0[30:21], 1'h0 };
  assign imm_s_type_o = { instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31:25], instr_rdata_i[11:7] };
  assign imm_s_type_o_t0 = { instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31:25], instr_rdata_i_t0[11:7] };
  assign imm_u_type_o = { instr_rdata_i[31:12], 12'h000 };
  assign imm_u_type_o_t0 = { instr_rdata_i_t0[31:12], 12'h000 };
  assign rf_raddr_a_o = instr_rdata_i[19:15];
  assign rf_raddr_a_o_t0 = instr_rdata_i_t0[19:15];
  assign rf_raddr_b_o = instr_rdata_i[24:20];
  assign rf_raddr_b_o_t0 = instr_rdata_i_t0[24:20];
  assign rf_waddr_o = instr_rdata_i[11:7];
  assign rf_waddr_o_t0 = instr_rdata_i_t0[11:7];
  assign zimm_rs1_type_o = { 27'h0000000, instr_rdata_i[19:15] };
  assign zimm_rs1_type_o_t0 = { 27'h0000000, instr_rdata_i_t0[19:15] };
endmodule

module paramodb14a8c3636c7c0bb82862600beccd3d8da4d4a94auxy_noerr_tlul_adapter_sram (clk_i, rst_ni, tl_i, tl_o, en_ifetch_i, req_o, req_type_o, gnt_i, we_o, addr_o, wdata_o, wmask_o, intg_error_o, rdata_i, rvalid_i, rerror_i, addr_o_t0, tl_i_t0, tl_o_t0, en_ifetch_i_t0, gnt_i_t0
, intg_error_o_t0, rdata_i_t0, req_o_t0, req_type_o_t0, rerror_i_t0, rvalid_i_t0, wdata_o_t0, we_o_t0, wmask_o_t0);
  wire [31:0] _0000_;
  wire [31:0] _0001_;
  wire [31:0] _0002_;
  wire [31:0] _0003_;
  wire [31:0] _0004_;
  wire [31:0] _0005_;
  wire [31:0] _0006_;
  wire [31:0] _0007_;
  wire [31:0] _0008_;
  wire [31:0] _0009_;
  wire [31:0] _0010_;
  wire [31:0] _0011_;
  wire [31:0] _0012_;
  wire [31:0] _0013_;
  wire [31:0] _0014_;
  wire [31:0] _0015_;
  wire [31:0] _0016_;
  wire [31:0] _0017_;
  wire [31:0] _0018_;
  wire [31:0] _0019_;
  wire [31:0] _0020_;
  wire [31:0] _0021_;
  wire _0022_;
  wire _0023_;
  wire _0024_;
  wire _0025_;
  wire _0026_;
  wire _0027_;
  wire [31:0] _0028_;
  wire [31:0] _0029_;
  wire [31:0] _0030_;
  wire [31:0] _0031_;
  wire [31:0] _0032_;
  wire [31:0] _0033_;
  wire [31:0] _0034_;
  wire [31:0] _0035_;
  wire [31:0] _0036_;
  wire [31:0] _0037_;
  wire [31:0] _0038_;
  wire [31:0] _0039_;
  wire [31:0] _0040_;
  wire [31:0] _0041_;
  wire [31:0] _0042_;
  wire [31:0] _0043_;
  wire [31:0] _0044_;
  wire [31:0] _0045_;
  wire [31:0] _0046_;
  wire [31:0] _0047_;
  wire [31:0] _0048_;
  wire [31:0] _0049_;
  wire [31:0] _0050_;
  wire [31:0] _0051_;
  wire [31:0] _0052_;
  wire [31:0] _0053_;
  wire [31:0] _0054_;
  wire [31:0] _0055_;
  wire [31:0] _0056_;
  wire [31:0] _0057_;
  wire [31:0] _0058_;
  wire [31:0] _0059_;
  wire [31:0] _0060_;
  wire [31:0] _0061_;
  wire [31:0] _0062_;
  wire [31:0] _0063_;
  wire [31:0] _0064_;
  wire [31:0] _0065_;
  wire [31:0] _0066_;
  wire [31:0] _0067_;
  wire [31:0] _0068_;
  wire [31:0] _0069_;
  wire [31:0] _0070_;
  wire [31:0] _0071_;
  wire _0072_;
  wire _0073_;
  wire _0074_;
  wire _0075_;
  wire [31:0] _0076_;
  wire [1:0] _0077_;
  wire [2:0] _0078_;
  wire [32:0] _0079_;
  wire [32:0] _0080_;
  wire [32:0] _0081_;
  wire [32:0] _0082_;
  wire [31:0] _0083_;
  wire [31:0] _0084_;
  wire [31:0] _0085_;
  wire [31:0] _0086_;
  wire [31:0] _0087_;
  wire [31:0] _0088_;
  wire [31:0] _0089_;
  wire [31:0] _0090_;
  wire [31:0] _0091_;
  wire [31:0] _0092_;
  wire [31:0] _0093_;
  wire [31:0] _0094_;
  wire [31:0] _0095_;
  wire [31:0] _0096_;
  wire [31:0] _0097_;
  wire [31:0] _0098_;
  wire [31:0] _0099_;
  wire [31:0] _0100_;
  wire [31:0] _0101_;
  wire [31:0] _0102_;
  wire _0103_;
  wire _0104_;
  wire [31:0] _0105_;
  wire _0106_;
  wire [1:0] _0107_;
  wire [2:0] _0108_;
  wire [6:0] _0109_;
  wire [31:0] _0110_;
  wire [7:0] _0111_;
  wire [1:0] _0112_;
  wire [17:0] _0113_;
  wire [7:0] _0114_;
  wire [7:0] _0115_;
  wire [7:0] _0116_;
  wire [7:0] _0117_;
  wire [1:0] _0118_;
  wire _0119_;
  wire _0120_;
  wire [32:0] _0121_;
  wire [32:0] _0122_;
  wire [32:0] _0123_;
  wire [32:0] _0124_;
  wire [32:0] _0125_;
  wire [32:0] _0126_;
  wire [32:0] _0127_;
  wire [32:0] _0128_;
  wire _0129_;
  wire _0130_;
  wire _0131_;
  wire _0132_;
  wire _0133_;
  wire _0134_;
  wire _0135_;
  wire _0136_;
  wire [31:0] _0137_;
  wire [31:0] _0138_;
  wire [31:0] _0139_;
  wire [31:0] _0140_;
  wire [31:0] _0141_;
  wire [31:0] _0142_;
  wire [31:0] _0143_;
  wire [31:0] _0144_;
  wire [31:0] _0145_;
  wire [31:0] _0146_;
  wire [31:0] _0147_;
  wire [31:0] _0148_;
  wire [31:0] _0149_;
  wire [31:0] _0150_;
  wire [31:0] _0151_;
  wire [31:0] _0152_;
  wire [31:0] _0153_;
  wire [31:0] _0154_;
  wire [31:0] _0155_;
  wire [31:0] _0156_;
  wire [31:0] _0157_;
  wire [31:0] _0158_;
  wire [31:0] _0159_;
  wire [31:0] _0160_;
  wire [31:0] _0161_;
  wire [31:0] _0162_;
  wire [31:0] _0163_;
  wire [31:0] _0164_;
  wire [31:0] _0165_;
  wire [31:0] _0166_;
  wire [31:0] _0167_;
  wire [31:0] _0168_;
  wire [31:0] _0169_;
  wire [31:0] _0170_;
  wire [31:0] _0171_;
  wire [31:0] _0172_;
  wire [31:0] _0173_;
  wire [31:0] _0174_;
  wire [31:0] _0175_;
  wire [31:0] _0176_;
  wire [31:0] _0177_;
  wire [31:0] _0178_;
  wire [31:0] _0179_;
  wire [31:0] _0180_;
  wire [31:0] _0181_;
  wire [31:0] _0182_;
  wire [31:0] _0183_;
  wire [31:0] _0184_;
  wire [31:0] _0185_;
  wire [31:0] _0186_;
  wire [31:0] _0187_;
  wire [31:0] _0188_;
  wire [31:0] _0189_;
  wire [31:0] _0190_;
  wire [31:0] _0191_;
  wire [31:0] _0192_;
  wire [31:0] _0193_;
  wire [31:0] _0194_;
  wire [31:0] _0195_;
  wire [31:0] _0196_;
  wire [31:0] _0197_;
  wire [31:0] _0198_;
  wire [31:0] _0199_;
  wire [31:0] _0200_;
  wire [31:0] _0201_;
  wire _0202_;
  wire _0203_;
  wire _0204_;
  wire _0205_;
  wire _0206_;
  wire _0207_;
  wire _0208_;
  wire _0209_;
  wire _0210_;
  wire _0211_;
  wire _0212_;
  wire _0213_;
  wire _0214_;
  wire _0215_;
  wire _0216_;
  wire _0217_;
  wire _0218_;
  wire _0219_;
  wire _0220_;
  wire _0221_;
  wire _0222_;
  wire _0223_;
  wire _0224_;
  wire _0225_;
  wire _0226_;
  wire _0227_;
  wire _0228_;
  wire [31:0] _0229_;
  wire [31:0] _0230_;
  wire [31:0] _0231_;
  wire _0232_;
  wire _0233_;
  wire _0234_;
  wire [1:0] _0235_;
  wire [1:0] _0236_;
  wire _0237_;
  wire _0238_;
  wire _0239_;
  wire _0240_;
  wire _0241_;
  wire _0242_;
  wire _0243_;
  wire _0244_;
  wire _0245_;
  wire _0246_;
  wire _0247_;
  wire _0248_;
  wire _0249_;
  wire _0250_;
  wire _0251_;
  wire _0252_;
  wire _0253_;
  wire _0254_;
  wire _0255_;
  wire _0256_;
  wire _0257_;
  wire _0258_;
  wire _0259_;
  wire _0260_;
  wire [2:0] _0261_;
  wire [2:0] _0262_;
  wire [32:0] _0263_;
  wire [32:0] _0264_;
  wire [32:0] _0265_;
  wire [32:0] _0266_;
  wire [31:0] _0267_;
  wire [31:0] _0268_;
  wire [31:0] _0269_;
  wire [31:0] _0270_;
  wire [31:0] _0271_;
  wire [31:0] _0272_;
  wire [31:0] _0273_;
  wire [31:0] _0274_;
  wire [31:0] _0275_;
  wire [31:0] _0276_;
  wire [31:0] _0277_;
  wire [31:0] _0278_;
  wire [31:0] _0279_;
  wire [31:0] _0280_;
  wire [31:0] _0281_;
  wire [31:0] _0282_;
  wire [31:0] _0283_;
  wire [31:0] _0284_;
  wire [31:0] _0285_;
  wire [31:0] _0286_;
  wire [31:0] _0287_;
  wire [31:0] _0288_;
  wire [31:0] _0289_;
  wire [31:0] _0290_;
  wire [31:0] _0291_;
  wire [31:0] _0292_;
  wire [31:0] _0293_;
  wire [31:0] _0294_;
  wire [31:0] _0295_;
  wire [31:0] _0296_;
  wire _0297_;
  wire _0298_;
  wire _0299_;
  wire [31:0] _0300_;
  wire [31:0] _0301_;
  wire [31:0] _0302_;
  wire [31:0] _0303_;
  wire [31:0] _0304_;
  wire _0305_;
  wire _0306_;
  wire _0307_;
  wire _0308_;
  wire _0309_;
  wire _0310_;
  wire _0311_;
  wire _0312_;
  wire _0313_;
  wire _0314_;
  wire _0315_;
  wire [1:0] _0316_;
  wire [2:0] _0317_;
  wire [2:0] _0318_;
  wire [2:0] _0319_;
  wire [6:0] _0320_;
  wire [6:0] _0321_;
  wire [6:0] _0322_;
  wire [31:0] _0323_;
  wire [31:0] _0324_;
  wire [31:0] _0325_;
  wire [7:0] _0326_;
  wire [7:0] _0327_;
  wire [7:0] _0328_;
  wire [1:0] _0329_;
  wire [1:0] _0330_;
  wire [1:0] _0331_;
  wire [17:0] _0332_;
  wire [17:0] _0333_;
  wire [17:0] _0334_;
  wire [7:0] _0335_;
  wire [7:0] _0336_;
  wire [7:0] _0337_;
  wire [7:0] _0338_;
  wire [7:0] _0339_;
  wire [7:0] _0340_;
  wire [7:0] _0341_;
  wire [7:0] _0342_;
  wire [7:0] _0343_;
  wire [7:0] _0344_;
  wire [7:0] _0345_;
  wire [7:0] _0346_;
  wire [1:0] _0347_;
  wire [1:0] _0348_;
  wire [1:0] _0349_;
  wire _0350_;
  wire _0351_;
  wire [31:0] _0352_;
  wire [31:0] _0353_;
  wire [31:0] _0354_;
  wire [31:0] _0355_;
  wire [31:0] _0356_;
  wire [31:0] _0357_;
  wire [31:0] _0358_;
  wire [31:0] _0359_;
  wire [31:0] _0360_;
  wire [31:0] _0361_;
  wire [31:0] _0362_;
  wire [31:0] _0363_;
  wire [31:0] _0364_;
  wire [31:0] _0365_;
  wire [31:0] _0366_;
  wire [31:0] _0367_;
  wire [31:0] _0368_;
  wire [31:0] _0369_;
  wire [31:0] _0370_;
  wire [31:0] _0371_;
  wire [31:0] _0372_;
  wire [31:0] _0373_;
  wire [31:0] _0374_;
  wire _0375_;
  wire _0376_;
  wire _0377_;
  wire _0378_;
  wire _0379_;
  wire _0380_;
  wire _0381_;
  wire _0382_;
  wire _0383_;
  wire [31:0] _0384_;
  wire _0385_;
  wire _0386_;
  wire _0387_;
  wire _0388_;
  wire _0389_;
  wire _0390_;
  wire _0391_;
  wire _0392_;
  wire _0393_;
  wire [32:0] _0394_;
  wire [32:0] _0395_;
  wire [32:0] _0396_;
  wire [32:0] _0397_;
  wire [31:0] _0398_;
  wire [31:0] _0399_;
  wire [31:0] _0400_;
  wire [31:0] _0401_;
  wire [31:0] _0402_;
  wire [31:0] _0403_;
  wire [31:0] _0404_;
  wire [31:0] _0405_;
  wire [31:0] _0406_;
  wire [31:0] _0407_;
  wire _0408_;
  wire [31:0] _0409_;
  wire [31:0] _0410_;
  wire [31:0] _0411_;
  wire [31:0] _0412_;
  wire _0413_;
  wire _0414_;
  wire _0415_;
  wire _0416_;
  wire _0417_;
  wire [2:0] _0418_;
  wire [2:0] _0419_;
  wire [2:0] _0420_;
  wire [6:0] _0421_;
  wire [6:0] _0422_;
  wire [6:0] _0423_;
  wire [31:0] _0424_;
  wire [31:0] _0425_;
  wire [31:0] _0426_;
  wire [7:0] _0427_;
  wire [7:0] _0428_;
  wire [7:0] _0429_;
  wire [1:0] _0430_;
  wire [1:0] _0431_;
  wire [1:0] _0432_;
  wire [17:0] _0433_;
  wire [17:0] _0434_;
  wire [17:0] _0435_;
  wire [7:0] _0436_;
  wire [7:0] _0437_;
  wire [7:0] _0438_;
  wire [7:0] _0439_;
  wire [7:0] _0440_;
  wire [7:0] _0441_;
  wire [7:0] _0442_;
  wire [7:0] _0443_;
  wire [7:0] _0444_;
  wire [7:0] _0445_;
  wire [7:0] _0446_;
  wire [7:0] _0447_;
  wire [1:0] _0448_;
  wire [1:0] _0449_;
  wire [1:0] _0450_;
  wire _0451_;
  wire [31:0] _0452_;
  wire [31:0] _0453_;
  wire [31:0] _0454_;
  wire [32:0] _0455_;
  wire [32:0] _0456_;
  wire [32:0] _0457_;
  wire [32:0] _0458_;
  wire [31:0] _0459_;
  wire [31:0] _0460_;
  wire _0461_;
  wire [6:0] _0462_;
  wire _0463_;
  wire _0464_;
  wire [31:0] _0465_;
  wire [31:0] _0466_;
  wire [31:0] _0467_;
  wire [31:0] _0468_;
  wire [31:0] _0469_;
  wire [31:0] _0470_;
  wire [31:0] _0471_;
  wire [31:0] _0472_;
  wire [31:0] _0473_;
  wire [31:0] _0474_;
  wire [31:0] _0475_;
  wire [31:0] _0476_;
  wire [31:0] _0477_;
  wire [31:0] _0478_;
  wire [31:0] _0479_;
  wire _0480_;
  wire _0481_;
  wire _0482_;
  wire _0483_;
  wire _0484_;
  wire _0485_;
  wire _0486_;
  wire _0487_;
  wire _0488_;
  wire _0489_;
  wire _0490_;
  wire _0491_;
  wire _0492_;
  wire _0493_;
  wire _0494_;
  wire _0495_;
  wire _0496_;
  wire _0497_;
  wire _0498_;
  wire _0499_;
  wire _0500_;
  wire [32:0] _0501_;
  wire [32:0] _0502_;
  wire [32:0] _0503_;
  wire [32:0] _0504_;
  wire [32:0] _0505_;
  wire [32:0] _0506_;
  wire [32:0] _0507_;
  wire [32:0] _0508_;
  wire [31:0] _0509_;
  wire [31:0] _0510_;
  wire [31:0] _0511_;
  wire [31:0] _0512_;
  wire _0513_;
  wire [31:0] _0514_;
  wire [31:0] _0515_;
  wire [31:0] _0516_;
  wire [31:0] _0517_;
  wire [31:0] _0518_;
  wire [31:0] _0519_;
  wire [31:0] _0520_;
  wire [31:0] _0521_;
  wire [31:0] _0522_;
  wire [31:0] _0523_;
  wire [31:0] _0524_;
  wire [31:0] _0525_;
  wire [31:0] _0526_;
  wire [31:0] _0527_;
  wire [31:0] _0528_;
  wire [31:0] _0529_;
  wire _0530_;
  wire _0531_;
  wire _0532_;
  wire [7:0] _0533_;
  wire [7:0] _0534_;
  wire [7:0] _0535_;
  wire [7:0] _0536_;
  wire [7:0] _0537_;
  wire [7:0] _0538_;
  wire [7:0] _0539_;
  wire [7:0] _0540_;
  wire a_ack;
  wire a_ack_t0;
  output [17:0] addr_o;
  wire [17:0] addr_o;
  output [17:0] addr_o_t0;
  wire [17:0] addr_o_t0;
  input clk_i;
  wire clk_i;
  wire d_ack;
  wire d_ack_t0;
  wire d_error;
  wire d_error_t0;
  wire d_valid;
  wire d_valid_t0;
  input [2:0] en_ifetch_i;
  wire [2:0] en_ifetch_i;
  input [2:0] en_ifetch_i_t0;
  wire [2:0] en_ifetch_i_t0;
  input gnt_i;
  wire gnt_i;
  input gnt_i_t0;
  wire gnt_i_t0;
  output intg_error_o;
  wire intg_error_o;
  output intg_error_o_t0;
  wire intg_error_o_t0;
  wire [31:0] rdata;
  input [31:0] rdata_i;
  wire [31:0] rdata_i;
  input [31:0] rdata_i_t0;
  wire [31:0] rdata_i_t0;
  wire [31:0] rdata_t0;
  wire [31:0] rdata_tlword;
  wire [31:0] rdata_tlword_t0;
  output req_o;
  wire req_o;
  output req_o_t0;
  wire req_o_t0;
  output [1:0] req_type_o;
  wire [1:0] req_type_o;
  output [1:0] req_type_o_t0;
  wire [1:0] req_type_o_t0;
  wire [12:0] reqfifo_rdata;
  wire [12:0] reqfifo_rdata_t0;
  wire reqfifo_rvalid;
  wire reqfifo_rvalid_t0;
  wire [12:0] reqfifo_wdata;
  wire [12:0] reqfifo_wdata_t0;
  wire reqfifo_wready;
  wire reqfifo_wready_t0;
  input [1:0] rerror_i;
  wire [1:0] rerror_i;
  input [1:0] rerror_i_t0;
  wire [1:0] rerror_i_t0;
  wire [31:0] rmask;
  wire [31:0] rmask_t0;
  wire [39:0] rspfifo_rdata;
  wire [39:0] rspfifo_rdata_t0;
  wire rspfifo_rready;
  wire rspfifo_rready_t0;
  wire rspfifo_rvalid;
  wire rspfifo_rvalid_t0;
  wire rspfifo_wready;
  wire rspfifo_wready_t0;
  wire rspfifo_wvalid;
  wire rspfifo_wvalid_t0;
  input rst_ni;
  wire rst_ni;
  input rvalid_i;
  wire rvalid_i;
  input rvalid_i_t0;
  wire rvalid_i_t0;
  wire sram_ack;
  wire sram_ack_t0;
  wire [4:0] sramreqfifo_rdata;
  wire [4:0] sramreqfifo_rdata_t0;
  wire sramreqfifo_wready;
  wire sramreqfifo_wready_t0;
  wire sramreqfifo_wvalid;
  wire sramreqfifo_wvalid_t0;
  wire [31:0] \sv2v_cast_35AE2$func$generated/sv2v_out.v:9139$93.$result ;
  wire [31:0] \sv2v_cast_35AE2$func$generated/sv2v_out.v:9139$93.$result_t0 ;
  wire [1:0] \sv2v_cast_4660A$func$generated/sv2v_out.v:9139$96.$result ;
  wire [1:0] \sv2v_cast_4660A$func$generated/sv2v_out.v:9139$96.$result_t0 ;
  wire [6:0] \sv2v_cast_8DC45$func$generated/sv2v_out.v:9139$90.$result ;
  wire [6:0] \sv2v_cast_8DC45$func$generated/sv2v_out.v:9139$90.$result_t0 ;
  wire [7:0] \sv2v_cast_964CB$func$generated/sv2v_out.v:9139$95.$result ;
  wire [7:0] \sv2v_cast_964CB$func$generated/sv2v_out.v:9139$95.$result_t0 ;
  input [106:0] tl_i;
  wire [106:0] tl_i;
  input [106:0] tl_i_t0;
  wire [106:0] tl_i_t0;
  output [65:0] tl_o;
  wire [65:0] tl_o;
  output [65:0] tl_o_t0;
  wire [65:0] tl_o_t0;
  wire [65:0] tl_out;
  wire [65:0] tl_out_t0;
  output [31:0] wdata_o;
  wire [31:0] wdata_o;
  output [31:0] wdata_o_t0;
  wire [31:0] wdata_o_t0;
  output we_o;
  wire we_o;
  output we_o_t0;
  wire we_o_t0;
  output [31:0] wmask_o;
  wire [31:0] wmask_o;
  output [31:0] wmask_o_t0;
  wire [31:0] wmask_o_t0;
  assign _0016_ = { 26'h0000000, sramreqfifo_rdata[0], 5'h00 } + 32'd8;
  assign _0018_ = { 26'h0000000, sramreqfifo_rdata[0], 5'h00 } + 32'd16;
  assign _0020_ = { 26'h0000000, sramreqfifo_rdata[0], 5'h00 } + 32'd24;
  assign _0028_ = 8'hff & { 24'h000000, tl_i[54], tl_i[54], tl_i[54], tl_i[54], tl_i[54], tl_i[54], tl_i[54], tl_i[54] };
  assign _0030_ = 8'hff & { 24'h000000, _0533_ };
  assign _0032_ = 8'hff & { 24'h000000, tl_i[55], tl_i[55], tl_i[55], tl_i[55], tl_i[55], tl_i[55], tl_i[55], tl_i[55] };
  assign _0034_ = _0028_ & 32'd4294902015;
  assign _0036_ = 8'hff & { 24'h000000, _0535_ };
  assign _0038_ = _0030_ & 32'd4294902015;
  assign _0040_ = 8'hff & { 24'h000000, tl_i[56], tl_i[56], tl_i[56], tl_i[56], tl_i[56], tl_i[56], tl_i[56], tl_i[56] };
  assign _0042_ = _0514_ & 32'd4278255615;
  assign _0044_ = 8'hff & { 24'h000000, _0537_ };
  assign _0046_ = _0516_ & 32'd4278255615;
  assign _0048_ = 8'hff & { 24'h000000, tl_i[57], tl_i[57], tl_i[57], tl_i[57], tl_i[57], tl_i[57], tl_i[57], tl_i[57] };
  assign _0050_ = _0518_ & 32'd16777215;
  assign _0052_ = 8'hff & { 24'h000000, _0539_ };
  assign _0054_ = _0520_ & 32'd16777215;
  assign _0056_ = 8'hff & { 24'h000000, sramreqfifo_rdata[1], sramreqfifo_rdata[1], sramreqfifo_rdata[1], sramreqfifo_rdata[1], sramreqfifo_rdata[1], sramreqfifo_rdata[1], sramreqfifo_rdata[1], sramreqfifo_rdata[1] };
  assign _0060_ = 8'hff & { 24'h000000, sramreqfifo_rdata[2], sramreqfifo_rdata[2], sramreqfifo_rdata[2], sramreqfifo_rdata[2], sramreqfifo_rdata[2], sramreqfifo_rdata[2], sramreqfifo_rdata[2], sramreqfifo_rdata[2] };
  assign _0062_ = _0524_ & _0510_;
  assign _0064_ = 8'hff & { 24'h000000, sramreqfifo_rdata[3], sramreqfifo_rdata[3], sramreqfifo_rdata[3], sramreqfifo_rdata[3], sramreqfifo_rdata[3], sramreqfifo_rdata[3], sramreqfifo_rdata[3], sramreqfifo_rdata[3] };
  assign _0066_ = _0526_ & _0511_;
  assign _0068_ = 8'hff & { 24'h000000, sramreqfifo_rdata[4], sramreqfifo_rdata[4], sramreqfifo_rdata[4], sramreqfifo_rdata[4], sramreqfifo_rdata[4], sramreqfifo_rdata[4], sramreqfifo_rdata[4], sramreqfifo_rdata[4] };
  assign _0070_ = _0528_ & _0512_;
  assign a_ack = tl_i[106] & tl_o[0];
  assign d_ack = tl_o[65] & tl_i[0];
  assign sram_ack = req_o & gnt_i;
  assign _0072_ = gnt_i & reqfifo_wready;
  assign tl_out[0] = _0072_ & sramreqfifo_wready;
  assign req_o = tl_i[106] & reqfifo_wready;
  assign we_o = tl_i[106] & _0496_;
  assign sramreqfifo_wvalid = sram_ack & _0513_;
  assign rspfifo_wvalid = rvalid_i & reqfifo_rvalid;
  assign rdata = rdata_i & rmask;
  assign _0074_ = _0480_ & _0104_;
  assign _0076_ = ~ { 26'h0000000, sramreqfifo_rdata_t0[0], 5'h00 };
  assign _0137_ = { 26'h0000000, sramreqfifo_rdata[0], 5'h00 } & _0076_;
  assign _0465_ = _0137_ + 32'd8;
  assign _0467_ = _0137_ + 32'd16;
  assign _0469_ = _0137_ + 32'd24;
  assign _0352_ = { 26'h0000000, sramreqfifo_rdata[0], 5'h00 } | { 26'h0000000, sramreqfifo_rdata_t0[0], 5'h00 };
  assign _0466_ = _0352_ + 32'd8;
  assign _0468_ = _0352_ + 32'd16;
  assign _0470_ = _0352_ + 32'd24;
  assign _0452_ = _0465_ ^ _0466_;
  assign _0453_ = _0467_ ^ _0468_;
  assign _0454_ = _0469_ ^ _0470_;
  assign _0017_ = _0452_ | { 26'h0000000, sramreqfifo_rdata_t0[0], 5'h00 };
  assign _0019_ = _0453_ | { 26'h0000000, sramreqfifo_rdata_t0[0], 5'h00 };
  assign _0021_ = _0454_ | { 26'h0000000, sramreqfifo_rdata_t0[0], 5'h00 };
  assign _0138_ = 32'd0 & { 24'h000000, tl_i[54], tl_i[54], tl_i[54], tl_i[54], tl_i[54], tl_i[54], tl_i[54], tl_i[54] };
  assign _0141_ = 32'd0 & { 24'h000000, _0533_ };
  assign _0144_ = 32'd0 & { 24'h000000, tl_i[55], tl_i[55], tl_i[55], tl_i[55], tl_i[55], tl_i[55], tl_i[55], tl_i[55] };
  assign _0147_ = _0029_ & 32'd4294902015;
  assign _0150_ = 32'd0 & { 24'h000000, _0535_ };
  assign _0153_ = _0031_ & 32'd4294902015;
  assign _0156_ = 32'd0 & { 24'h000000, tl_i[56], tl_i[56], tl_i[56], tl_i[56], tl_i[56], tl_i[56], tl_i[56], tl_i[56] };
  assign _0159_ = _0515_ & 32'd4278255615;
  assign _0162_ = 32'd0 & { 24'h000000, _0537_ };
  assign _0165_ = _0517_ & 32'd4278255615;
  assign _0168_ = 32'd0 & { 24'h000000, tl_i[57], tl_i[57], tl_i[57], tl_i[57], tl_i[57], tl_i[57], tl_i[57], tl_i[57] };
  assign _0171_ = _0519_ & 32'd16777215;
  assign _0174_ = 32'd0 & { 24'h000000, _0539_ };
  assign _0177_ = _0521_ & 32'd16777215;
  assign _0180_ = 32'd0 & { 24'h000000, sramreqfifo_rdata[1], sramreqfifo_rdata[1], sramreqfifo_rdata[1], sramreqfifo_rdata[1], sramreqfifo_rdata[1], sramreqfifo_rdata[1], sramreqfifo_rdata[1], sramreqfifo_rdata[1] };
  assign _0058_ = 32'd0 & _0509_;
  assign _0184_ = 32'd0 & { 24'h000000, sramreqfifo_rdata[2], sramreqfifo_rdata[2], sramreqfifo_rdata[2], sramreqfifo_rdata[2], sramreqfifo_rdata[2], sramreqfifo_rdata[2], sramreqfifo_rdata[2], sramreqfifo_rdata[2] };
  assign _0187_ = _0525_ & _0510_;
  assign _0190_ = 32'd0 & { 24'h000000, sramreqfifo_rdata[3], sramreqfifo_rdata[3], sramreqfifo_rdata[3], sramreqfifo_rdata[3], sramreqfifo_rdata[3], sramreqfifo_rdata[3], sramreqfifo_rdata[3], sramreqfifo_rdata[3] };
  assign _0193_ = _0527_ & _0511_;
  assign _0196_ = 32'd0 & { 24'h000000, sramreqfifo_rdata[4], sramreqfifo_rdata[4], sramreqfifo_rdata[4], sramreqfifo_rdata[4], sramreqfifo_rdata[4], sramreqfifo_rdata[4], sramreqfifo_rdata[4], sramreqfifo_rdata[4] };
  assign _0199_ = _0529_ & _0512_;
  assign _0202_ = tl_i_t0[106] & tl_o[0];
  assign _0205_ = tl_o_t0[65] & tl_i[0];
  assign _0208_ = req_o_t0 & gnt_i;
  assign _0211_ = gnt_i_t0 & reqfifo_wready;
  assign _0214_ = _0073_ & sramreqfifo_wready;
  assign _0217_ = tl_i_t0[106] & reqfifo_wready;
  assign _0220_ = tl_i_t0[106] & _0496_;
  assign _0223_ = sram_ack_t0 & _0513_;
  assign _0226_ = rvalid_i_t0 & reqfifo_rvalid;
  assign _0229_ = rdata_i_t0 & rmask;
  assign _0232_ = _0481_ & _0104_;
  assign _0139_ = { 24'h000000, tl_i_t0[54], tl_i_t0[54], tl_i_t0[54], tl_i_t0[54], tl_i_t0[54], tl_i_t0[54], tl_i_t0[54], tl_i_t0[54] } & 32'd255;
  assign _0142_ = { 24'h000000, _0534_ } & 32'd255;
  assign _0145_ = { 24'h000000, tl_i_t0[55], tl_i_t0[55], tl_i_t0[55], tl_i_t0[55], tl_i_t0[55], tl_i_t0[55], tl_i_t0[55], tl_i_t0[55] } & 32'd255;
  assign _0148_ = 32'd0 & _0028_;
  assign _0151_ = { 24'h000000, _0536_ } & 32'd255;
  assign _0154_ = 32'd0 & _0030_;
  assign _0157_ = { 24'h000000, tl_i_t0[56], tl_i_t0[56], tl_i_t0[56], tl_i_t0[56], tl_i_t0[56], tl_i_t0[56], tl_i_t0[56], tl_i_t0[56] } & 32'd255;
  assign _0160_ = 32'd0 & _0514_;
  assign _0163_ = { 24'h000000, _0538_ } & 32'd255;
  assign _0166_ = 32'd0 & _0516_;
  assign _0169_ = { 24'h000000, tl_i_t0[57], tl_i_t0[57], tl_i_t0[57], tl_i_t0[57], tl_i_t0[57], tl_i_t0[57], tl_i_t0[57], tl_i_t0[57] } & 32'd255;
  assign _0172_ = 32'd0 & _0518_;
  assign _0175_ = { 24'h000000, _0540_ } & 32'd255;
  assign _0178_ = 32'd0 & _0520_;
  assign _0181_ = { 24'h000000, sramreqfifo_rdata_t0[1], sramreqfifo_rdata_t0[1], sramreqfifo_rdata_t0[1], sramreqfifo_rdata_t0[1], sramreqfifo_rdata_t0[1], sramreqfifo_rdata_t0[1], sramreqfifo_rdata_t0[1], sramreqfifo_rdata_t0[1] } & 32'd255;
  assign _0185_ = { 24'h000000, sramreqfifo_rdata_t0[2], sramreqfifo_rdata_t0[2], sramreqfifo_rdata_t0[2], sramreqfifo_rdata_t0[2], sramreqfifo_rdata_t0[2], sramreqfifo_rdata_t0[2], sramreqfifo_rdata_t0[2], sramreqfifo_rdata_t0[2] } & 32'd255;
  assign _0188_ = _0011_ & _0524_;
  assign _0191_ = { 24'h000000, sramreqfifo_rdata_t0[3], sramreqfifo_rdata_t0[3], sramreqfifo_rdata_t0[3], sramreqfifo_rdata_t0[3], sramreqfifo_rdata_t0[3], sramreqfifo_rdata_t0[3], sramreqfifo_rdata_t0[3], sramreqfifo_rdata_t0[3] } & 32'd255;
  assign _0194_ = _0013_ & _0526_;
  assign _0197_ = { 24'h000000, sramreqfifo_rdata_t0[4], sramreqfifo_rdata_t0[4], sramreqfifo_rdata_t0[4], sramreqfifo_rdata_t0[4], sramreqfifo_rdata_t0[4], sramreqfifo_rdata_t0[4], sramreqfifo_rdata_t0[4], sramreqfifo_rdata_t0[4] } & 32'd255;
  assign _0200_ = _0015_ & _0528_;
  assign _0203_ = tl_o_t0[0] & tl_i[106];
  assign _0206_ = tl_i_t0[0] & tl_o[65];
  assign _0209_ = gnt_i_t0 & req_o;
  assign _0212_ = reqfifo_wready_t0 & gnt_i;
  assign _0215_ = sramreqfifo_wready_t0 & _0072_;
  assign _0218_ = reqfifo_wready_t0 & tl_i[106];
  assign _0221_ = _0497_ & tl_i[106];
  assign _0224_ = we_o_t0 & sram_ack;
  assign _0227_ = reqfifo_rvalid_t0 & rvalid_i;
  assign _0230_ = rmask_t0 & rdata_i;
  assign _0233_ = reqfifo_rdata_t0[10] & _0480_;
  assign _0140_ = 32'd0 & { 24'h000000, tl_i_t0[54], tl_i_t0[54], tl_i_t0[54], tl_i_t0[54], tl_i_t0[54], tl_i_t0[54], tl_i_t0[54], tl_i_t0[54] };
  assign _0143_ = 32'd0 & { 24'h000000, _0534_ };
  assign _0146_ = 32'd0 & { 24'h000000, tl_i_t0[55], tl_i_t0[55], tl_i_t0[55], tl_i_t0[55], tl_i_t0[55], tl_i_t0[55], tl_i_t0[55], tl_i_t0[55] };
  assign _0149_ = _0029_ & 32'd0;
  assign _0152_ = 32'd0 & { 24'h000000, _0536_ };
  assign _0155_ = _0031_ & 32'd0;
  assign _0158_ = 32'd0 & { 24'h000000, tl_i_t0[56], tl_i_t0[56], tl_i_t0[56], tl_i_t0[56], tl_i_t0[56], tl_i_t0[56], tl_i_t0[56], tl_i_t0[56] };
  assign _0161_ = _0515_ & 32'd0;
  assign _0164_ = 32'd0 & { 24'h000000, _0538_ };
  assign _0167_ = _0517_ & 32'd0;
  assign _0170_ = 32'd0 & { 24'h000000, tl_i_t0[57], tl_i_t0[57], tl_i_t0[57], tl_i_t0[57], tl_i_t0[57], tl_i_t0[57], tl_i_t0[57], tl_i_t0[57] };
  assign _0173_ = _0519_ & 32'd0;
  assign _0176_ = 32'd0 & { 24'h000000, _0540_ };
  assign _0179_ = _0521_ & 32'd0;
  assign _0182_ = 32'd0 & { 24'h000000, sramreqfifo_rdata_t0[1], sramreqfifo_rdata_t0[1], sramreqfifo_rdata_t0[1], sramreqfifo_rdata_t0[1], sramreqfifo_rdata_t0[1], sramreqfifo_rdata_t0[1], sramreqfifo_rdata_t0[1], sramreqfifo_rdata_t0[1] };
  assign _0183_ = 32'd0 & _0009_;
  assign _0186_ = 32'd0 & { 24'h000000, sramreqfifo_rdata_t0[2], sramreqfifo_rdata_t0[2], sramreqfifo_rdata_t0[2], sramreqfifo_rdata_t0[2], sramreqfifo_rdata_t0[2], sramreqfifo_rdata_t0[2], sramreqfifo_rdata_t0[2], sramreqfifo_rdata_t0[2] };
  assign _0189_ = _0525_ & _0011_;
  assign _0192_ = 32'd0 & { 24'h000000, sramreqfifo_rdata_t0[3], sramreqfifo_rdata_t0[3], sramreqfifo_rdata_t0[3], sramreqfifo_rdata_t0[3], sramreqfifo_rdata_t0[3], sramreqfifo_rdata_t0[3], sramreqfifo_rdata_t0[3], sramreqfifo_rdata_t0[3] };
  assign _0195_ = _0527_ & _0013_;
  assign _0198_ = 32'd0 & { 24'h000000, sramreqfifo_rdata_t0[4], sramreqfifo_rdata_t0[4], sramreqfifo_rdata_t0[4], sramreqfifo_rdata_t0[4], sramreqfifo_rdata_t0[4], sramreqfifo_rdata_t0[4], sramreqfifo_rdata_t0[4], sramreqfifo_rdata_t0[4] };
  assign _0201_ = _0529_ & _0015_;
  assign _0204_ = tl_i_t0[106] & tl_o_t0[0];
  assign _0207_ = tl_o_t0[65] & tl_i_t0[0];
  assign _0210_ = req_o_t0 & gnt_i_t0;
  assign _0213_ = gnt_i_t0 & reqfifo_wready_t0;
  assign _0216_ = _0073_ & sramreqfifo_wready_t0;
  assign _0219_ = tl_i_t0[106] & reqfifo_wready_t0;
  assign _0222_ = tl_i_t0[106] & _0497_;
  assign _0225_ = sram_ack_t0 & we_o_t0;
  assign _0228_ = rvalid_i_t0 & reqfifo_rvalid_t0;
  assign _0231_ = rdata_i_t0 & rmask_t0;
  assign _0234_ = _0481_ & reqfifo_rdata_t0[10];
  assign _0353_ = _0138_ | _0139_;
  assign _0354_ = _0141_ | _0142_;
  assign _0355_ = _0144_ | _0145_;
  assign _0356_ = _0147_ | _0148_;
  assign _0357_ = _0150_ | _0151_;
  assign _0358_ = _0153_ | _0154_;
  assign _0359_ = _0156_ | _0157_;
  assign _0360_ = _0159_ | _0160_;
  assign _0361_ = _0162_ | _0163_;
  assign _0362_ = _0165_ | _0166_;
  assign _0363_ = _0168_ | _0169_;
  assign _0364_ = _0171_ | _0172_;
  assign _0365_ = _0174_ | _0175_;
  assign _0366_ = _0177_ | _0178_;
  assign _0367_ = _0180_ | _0181_;
  assign _0368_ = _0058_ | _0183_;
  assign _0369_ = _0184_ | _0185_;
  assign _0370_ = _0187_ | _0188_;
  assign _0371_ = _0190_ | _0191_;
  assign _0372_ = _0193_ | _0194_;
  assign _0373_ = _0196_ | _0197_;
  assign _0374_ = _0199_ | _0200_;
  assign _0375_ = _0202_ | _0203_;
  assign _0376_ = _0205_ | _0206_;
  assign _0377_ = _0208_ | _0209_;
  assign _0378_ = _0211_ | _0212_;
  assign _0379_ = _0214_ | _0215_;
  assign _0380_ = _0217_ | _0218_;
  assign _0381_ = _0220_ | _0221_;
  assign _0382_ = _0223_ | _0224_;
  assign _0383_ = _0226_ | _0227_;
  assign _0384_ = _0229_ | _0230_;
  assign _0385_ = _0232_ | _0233_;
  assign _0029_ = _0353_ | _0140_;
  assign _0031_ = _0354_ | _0143_;
  assign _0033_ = _0355_ | _0146_;
  assign _0035_ = _0356_ | _0149_;
  assign _0037_ = _0357_ | _0152_;
  assign _0039_ = _0358_ | _0155_;
  assign _0041_ = _0359_ | _0158_;
  assign _0043_ = _0360_ | _0161_;
  assign _0045_ = _0361_ | _0164_;
  assign _0047_ = _0362_ | _0167_;
  assign _0049_ = _0363_ | _0170_;
  assign _0051_ = _0364_ | _0173_;
  assign _0053_ = _0365_ | _0176_;
  assign _0055_ = _0366_ | _0179_;
  assign _0057_ = _0367_ | _0182_;
  assign _0059_ = _0368_ | _0183_;
  assign _0061_ = _0369_ | _0186_;
  assign _0063_ = _0370_ | _0189_;
  assign _0065_ = _0371_ | _0192_;
  assign _0067_ = _0372_ | _0195_;
  assign _0069_ = _0373_ | _0198_;
  assign _0071_ = _0374_ | _0201_;
  assign a_ack_t0 = _0375_ | _0204_;
  assign d_ack_t0 = _0376_ | _0207_;
  assign sram_ack_t0 = _0377_ | _0210_;
  assign _0073_ = _0378_ | _0213_;
  assign tl_out_t0[0] = _0379_ | _0216_;
  assign req_o_t0 = _0380_ | _0219_;
  assign we_o_t0 = _0381_ | _0222_;
  assign sramreqfifo_wvalid_t0 = _0382_ | _0225_;
  assign rspfifo_wvalid_t0 = _0383_ | _0228_;
  assign rdata_t0 = _0384_ | _0231_;
  assign _0075_ = _0385_ | _0234_;
  assign _0129_ = | reqfifo_rdata_t0[12:11];
  assign _0130_ = | tl_i_t0[105:103];
  assign _0077_ = ~ reqfifo_rdata_t0[12:11];
  assign _0078_ = ~ tl_i_t0[105:103];
  assign _0235_ = reqfifo_rdata[12:11] & _0077_;
  assign _0261_ = tl_i[105:103] & _0078_;
  assign _0236_ = 2'h1 & _0077_;
  assign _0262_ = 3'h4 & _0078_;
  assign _0463_ = _0235_ == _0236_;
  assign _0464_ = _0261_ == _0262_;
  assign _0481_ = _0463_ & _0129_;
  assign _0500_ = _0464_ & _0130_;
  assign _0237_ = d_valid_t0 & d_error;
  assign _0240_ = d_valid_t0 & _0498_;
  assign _0243_ = d_valid_t0 & rspfifo_rvalid;
  assign _0246_ = _0485_ & _0480_;
  assign _0249_ = tl_i_t0[54] & we_o;
  assign _0252_ = tl_i_t0[55] & we_o;
  assign _0255_ = tl_i_t0[56] & we_o;
  assign _0258_ = tl_i_t0[57] & we_o;
  assign _0238_ = d_error_t0 & d_valid;
  assign _0241_ = _0481_ & d_valid;
  assign _0244_ = rspfifo_rvalid_t0 & d_valid;
  assign _0247_ = _0481_ & _0484_;
  assign _0250_ = we_o_t0 & tl_i[54];
  assign _0253_ = we_o_t0 & tl_i[55];
  assign _0256_ = we_o_t0 & tl_i[56];
  assign _0259_ = we_o_t0 & tl_i[57];
  assign _0239_ = d_valid_t0 & d_error_t0;
  assign _0242_ = d_valid_t0 & _0481_;
  assign _0245_ = d_valid_t0 & rspfifo_rvalid_t0;
  assign _0248_ = _0485_ & _0481_;
  assign _0251_ = tl_i_t0[54] & we_o_t0;
  assign _0254_ = tl_i_t0[55] & we_o_t0;
  assign _0257_ = tl_i_t0[56] & we_o_t0;
  assign _0260_ = tl_i_t0[57] & we_o_t0;
  assign _0386_ = _0237_ | _0238_;
  assign _0387_ = _0240_ | _0241_;
  assign _0388_ = _0243_ | _0244_;
  assign _0389_ = _0246_ | _0247_;
  assign _0390_ = _0249_ | _0250_;
  assign _0391_ = _0252_ | _0253_;
  assign _0392_ = _0255_ | _0256_;
  assign _0393_ = _0258_ | _0259_;
  assign tl_out_t0[1] = _0386_ | _0239_;
  assign _0483_ = _0387_ | _0242_;
  assign _0485_ = _0388_ | _0245_;
  assign _0487_ = _0389_ | _0248_;
  assign _0489_ = _0390_ | _0251_;
  assign _0491_ = _0391_ | _0254_;
  assign _0493_ = _0392_ | _0257_;
  assign _0495_ = _0393_ | _0260_;
  assign _0131_ = | tl_i_t0[105:104];
  assign _0107_ = ~ tl_i_t0[105:104];
  assign _0316_ = tl_i[105:104] & _0107_;
  assign _0136_ = ! _0316_;
  assign _0497_ = _0136_ & _0131_;
  assign _0105_ = ~ { tl_i[106], tl_i[106], tl_i[106], tl_i[106], tl_i[106], tl_i[106], tl_i[106], tl_i[106], tl_i[106], tl_i[106], tl_i[106], tl_i[106], tl_i[106], tl_i[106], tl_i[106], tl_i[106], tl_i[106], tl_i[106], tl_i[106], tl_i[106], tl_i[106], tl_i[106], tl_i[106], tl_i[106], tl_i[106], tl_i[106], tl_i[106], tl_i[106], tl_i[106], tl_i[106], tl_i[106], tl_i[106] };
  assign _0106_ = ~ _0480_;
  assign _0104_ = ~ reqfifo_rdata[10];
  assign _0108_ = ~ { _0482_, _0482_, _0482_ };
  assign _0109_ = ~ { d_valid, d_valid, d_valid, d_valid, d_valid, d_valid, d_valid };
  assign _0110_ = ~ { _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_ };
  assign _0111_ = ~ { d_valid, d_valid, d_valid, d_valid, d_valid, d_valid, d_valid, d_valid };
  assign _0112_ = ~ { d_valid, d_valid };
  assign _0113_ = ~ { tl_i[106], tl_i[106], tl_i[106], tl_i[106], tl_i[106], tl_i[106], tl_i[106], tl_i[106], tl_i[106], tl_i[106], tl_i[106], tl_i[106], tl_i[106], tl_i[106], tl_i[106], tl_i[106], tl_i[106], tl_i[106] };
  assign _0114_ = ~ { _0488_, _0488_, _0488_, _0488_, _0488_, _0488_, _0488_, _0488_ };
  assign _0115_ = ~ { _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_ };
  assign _0116_ = ~ { _0492_, _0492_, _0492_, _0492_, _0492_, _0492_, _0492_, _0492_ };
  assign _0117_ = ~ { _0494_, _0494_, _0494_, _0494_, _0494_, _0494_, _0494_, _0494_ };
  assign _0118_ = ~ { _0499_, _0499_ };
  assign _0409_ = { tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106] } | _0105_;
  assign _0413_ = _0481_ | _0106_;
  assign _0417_ = reqfifo_rdata_t0[10] | _0104_;
  assign _0418_ = { _0483_, _0483_, _0483_ } | _0108_;
  assign _0421_ = { d_valid_t0, d_valid_t0, d_valid_t0, d_valid_t0, d_valid_t0, d_valid_t0, d_valid_t0 } | _0109_;
  assign _0424_ = { _0487_, _0487_, _0487_, _0487_, _0487_, _0487_, _0487_, _0487_, _0487_, _0487_, _0487_, _0487_, _0487_, _0487_, _0487_, _0487_, _0487_, _0487_, _0487_, _0487_, _0487_, _0487_, _0487_, _0487_, _0487_, _0487_, _0487_, _0487_, _0487_, _0487_, _0487_, _0487_ } | _0110_;
  assign _0427_ = { d_valid_t0, d_valid_t0, d_valid_t0, d_valid_t0, d_valid_t0, d_valid_t0, d_valid_t0, d_valid_t0 } | _0111_;
  assign _0430_ = { d_valid_t0, d_valid_t0 } | _0112_;
  assign _0433_ = { tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106] } | _0113_;
  assign _0436_ = { _0489_, _0489_, _0489_, _0489_, _0489_, _0489_, _0489_, _0489_ } | _0114_;
  assign _0439_ = { _0491_, _0491_, _0491_, _0491_, _0491_, _0491_, _0491_, _0491_ } | _0115_;
  assign _0442_ = { _0493_, _0493_, _0493_, _0493_, _0493_, _0493_, _0493_, _0493_ } | _0116_;
  assign _0445_ = { _0495_, _0495_, _0495_, _0495_, _0495_, _0495_, _0495_, _0495_ } | _0117_;
  assign _0448_ = { _0500_, _0500_ } | _0118_;
  assign _0410_ = { tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106] } | { tl_i[106], tl_i[106], tl_i[106], tl_i[106], tl_i[106], tl_i[106], tl_i[106], tl_i[106], tl_i[106], tl_i[106], tl_i[106], tl_i[106], tl_i[106], tl_i[106], tl_i[106], tl_i[106], tl_i[106], tl_i[106], tl_i[106], tl_i[106], tl_i[106], tl_i[106], tl_i[106], tl_i[106], tl_i[106], tl_i[106], tl_i[106], tl_i[106], tl_i[106], tl_i[106], tl_i[106], tl_i[106] };
  assign _0414_ = _0481_ | _0480_;
  assign _0416_ = reqfifo_rvalid_t0 | reqfifo_rvalid;
  assign _0419_ = { _0483_, _0483_, _0483_ } | { _0482_, _0482_, _0482_ };
  assign _0422_ = { d_valid_t0, d_valid_t0, d_valid_t0, d_valid_t0, d_valid_t0, d_valid_t0, d_valid_t0 } | { d_valid, d_valid, d_valid, d_valid, d_valid, d_valid, d_valid };
  assign _0425_ = { _0487_, _0487_, _0487_, _0487_, _0487_, _0487_, _0487_, _0487_, _0487_, _0487_, _0487_, _0487_, _0487_, _0487_, _0487_, _0487_, _0487_, _0487_, _0487_, _0487_, _0487_, _0487_, _0487_, _0487_, _0487_, _0487_, _0487_, _0487_, _0487_, _0487_, _0487_, _0487_ } | { _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_ };
  assign _0428_ = { d_valid_t0, d_valid_t0, d_valid_t0, d_valid_t0, d_valid_t0, d_valid_t0, d_valid_t0, d_valid_t0 } | { d_valid, d_valid, d_valid, d_valid, d_valid, d_valid, d_valid, d_valid };
  assign _0431_ = { d_valid_t0, d_valid_t0 } | { d_valid, d_valid };
  assign _0434_ = { tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106] } | { tl_i[106], tl_i[106], tl_i[106], tl_i[106], tl_i[106], tl_i[106], tl_i[106], tl_i[106], tl_i[106], tl_i[106], tl_i[106], tl_i[106], tl_i[106], tl_i[106], tl_i[106], tl_i[106], tl_i[106], tl_i[106] };
  assign _0437_ = { _0489_, _0489_, _0489_, _0489_, _0489_, _0489_, _0489_, _0489_ } | { _0488_, _0488_, _0488_, _0488_, _0488_, _0488_, _0488_, _0488_ };
  assign _0440_ = { _0491_, _0491_, _0491_, _0491_, _0491_, _0491_, _0491_, _0491_ } | { _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_ };
  assign _0443_ = { _0493_, _0493_, _0493_, _0493_, _0493_, _0493_, _0493_, _0493_ } | { _0492_, _0492_, _0492_, _0492_, _0492_, _0492_, _0492_, _0492_ };
  assign _0446_ = { _0495_, _0495_, _0495_, _0495_, _0495_, _0495_, _0495_, _0495_ } | { _0494_, _0494_, _0494_, _0494_, _0494_, _0494_, _0494_, _0494_ };
  assign _0449_ = { _0500_, _0500_ } | { _0499_, _0499_ };
  assign _0451_ = _0075_ | _0074_;
  assign _0300_ = 32'd0 & _0409_;
  assign _0305_ = reqfifo_rdata_t0[10] & _0413_;
  assign _0312_ = _0027_ & _0417_;
  assign _0317_ = 3'h0 & _0418_;
  assign _0320_ = 7'h00 & _0421_;
  assign _0323_ = 32'd0 & _0424_;
  assign _0326_ = 8'h00 & _0427_;
  assign _0329_ = 2'h0 & _0430_;
  assign _0332_ = 18'h00000 & _0433_;
  assign _0335_ = 8'h00 & _0436_;
  assign _0338_ = 8'h00 & _0439_;
  assign _0341_ = 8'h00 & _0442_;
  assign _0344_ = 8'h00 & _0445_;
  assign _0347_ = 2'h0 & _0448_;
  assign _0301_ = _0523_ & _0410_;
  assign _0303_ = _0522_ & _0410_;
  assign _0306_ = _0531_ & _0414_;
  assign _0308_ = _0023_ & _0416_;
  assign _0310_ = rspfifo_rvalid_t0 & _0414_;
  assign _0314_ = _0025_ & _0416_;
  assign _0318_ = 3'h0 & _0419_;
  assign _0321_ = rspfifo_rdata_t0[7:1] & _0422_;
  assign _0324_ = rspfifo_rdata_t0[39:8] & _0425_;
  assign _0327_ = reqfifo_rdata_t0[7:0] & _0428_;
  assign _0330_ = reqfifo_rdata_t0[9:8] & _0431_;
  assign _0333_ = tl_i_t0[77:60] & _0434_;
  assign _0336_ = tl_i_t0[29:22] & _0437_;
  assign _0339_ = tl_i_t0[37:30] & _0440_;
  assign _0342_ = tl_i_t0[45:38] & _0443_;
  assign _0345_ = tl_i_t0[53:46] & _0446_;
  assign _0348_ = 2'h0 & _0449_;
  assign _0350_ = d_ack_t0 & _0451_;
  assign _0411_ = _0300_ | _0301_;
  assign _0412_ = _0300_ | _0303_;
  assign _0415_ = _0305_ | _0306_;
  assign _0420_ = _0317_ | _0318_;
  assign _0423_ = _0320_ | _0321_;
  assign _0426_ = _0323_ | _0324_;
  assign _0429_ = _0326_ | _0327_;
  assign _0432_ = _0329_ | _0330_;
  assign _0435_ = _0332_ | _0333_;
  assign _0438_ = _0335_ | _0336_;
  assign _0441_ = _0338_ | _0339_;
  assign _0444_ = _0341_ | _0342_;
  assign _0447_ = _0344_ | _0345_;
  assign _0450_ = _0347_ | _0348_;
  assign _0461_ = reqfifo_rdata[10] ^ _0530_;
  assign _0462_ = 7'h7f ^ rspfifo_rdata[7:1];
  assign _0302_ = { tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106] } & _0459_;
  assign _0304_ = { tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106] } & _0460_;
  assign _0307_ = _0481_ & _0461_;
  assign _0309_ = reqfifo_rvalid_t0 & _0022_;
  assign _0311_ = _0481_ & _0119_;
  assign _0313_ = reqfifo_rdata_t0[10] & _0120_;
  assign _0315_ = reqfifo_rvalid_t0 & _0024_;
  assign _0319_ = { _0483_, _0483_, _0483_ } & 3'h1;
  assign _0322_ = { d_valid_t0, d_valid_t0, d_valid_t0, d_valid_t0, d_valid_t0, d_valid_t0, d_valid_t0 } & _0462_;
  assign _0325_ = { _0487_, _0487_, _0487_, _0487_, _0487_, _0487_, _0487_, _0487_, _0487_, _0487_, _0487_, _0487_, _0487_, _0487_, _0487_, _0487_, _0487_, _0487_, _0487_, _0487_, _0487_, _0487_, _0487_, _0487_, _0487_, _0487_, _0487_, _0487_, _0487_, _0487_, _0487_, _0487_ } & rspfifo_rdata[39:8];
  assign _0328_ = { d_valid_t0, d_valid_t0, d_valid_t0, d_valid_t0, d_valid_t0, d_valid_t0, d_valid_t0, d_valid_t0 } & reqfifo_rdata[7:0];
  assign _0331_ = { d_valid_t0, d_valid_t0 } & reqfifo_rdata[9:8];
  assign _0334_ = { tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106], tl_i_t0[106] } & tl_i[77:60];
  assign _0337_ = { _0489_, _0489_, _0489_, _0489_, _0489_, _0489_, _0489_, _0489_ } & tl_i[29:22];
  assign _0340_ = { _0491_, _0491_, _0491_, _0491_, _0491_, _0491_, _0491_, _0491_ } & tl_i[37:30];
  assign _0343_ = { _0493_, _0493_, _0493_, _0493_, _0493_, _0493_, _0493_, _0493_ } & tl_i[45:38];
  assign _0346_ = { _0495_, _0495_, _0495_, _0495_, _0495_, _0495_, _0495_, _0495_ } & tl_i[53:46];
  assign _0349_ = { _0500_, _0500_ } & 2'h1;
  assign _0351_ = _0075_ & d_ack;
  assign wdata_o_t0 = _0302_ | _0411_;
  assign wmask_o_t0 = _0304_ | _0412_;
  assign _0023_ = _0307_ | _0415_;
  assign d_error_t0 = _0309_ | _0308_;
  assign _0027_ = _0311_ | _0310_;
  assign _0025_ = _0313_ | _0312_;
  assign d_valid_t0 = _0315_ | _0314_;
  assign tl_out_t0[64:62] = _0319_ | _0420_;
  assign \sv2v_cast_8DC45$func$generated/sv2v_out.v:9139$90.$result_t0  = _0322_ | _0423_;
  assign \sv2v_cast_35AE2$func$generated/sv2v_out.v:9139$93.$result_t0  = _0325_ | _0426_;
  assign \sv2v_cast_964CB$func$generated/sv2v_out.v:9139$95.$result_t0  = _0328_ | _0429_;
  assign \sv2v_cast_4660A$func$generated/sv2v_out.v:9139$96.$result_t0  = _0331_ | _0432_;
  assign addr_o_t0 = _0334_ | _0435_;
  assign _0534_ = _0337_ | _0438_;
  assign _0536_ = _0340_ | _0441_;
  assign _0538_ = _0343_ | _0444_;
  assign _0540_ = _0346_ | _0447_;
  assign reqfifo_wdata_t0[12:11] = _0349_ | _0450_;
  assign rspfifo_rready_t0 = _0351_ | _0350_;
  assign _0079_ = ~ { 27'h0000000, sramreqfifo_rdata_t0[0], 5'h00 };
  assign _0080_ = ~ { 1'h0, _0017_ };
  assign _0081_ = ~ { 1'h0, _0019_ };
  assign _0082_ = ~ { 1'h0, _0021_ };
  assign _0263_ = { 27'h0000000, sramreqfifo_rdata[0], 5'h00 } & _0079_;
  assign _0264_ = { 1'h0, _0016_ } & _0080_;
  assign _0265_ = { 1'h0, _0018_ } & _0081_;
  assign _0266_ = { 1'h0, _0020_ } & _0082_;
  assign _0394_ = { 27'h0000000, sramreqfifo_rdata[0], 5'h00 } | { 27'h0000000, sramreqfifo_rdata_t0[0], 5'h00 };
  assign _0395_ = { 1'h0, _0016_ } | { 1'h0, _0017_ };
  assign _0396_ = { 1'h0, _0018_ } | { 1'h0, _0019_ };
  assign _0397_ = { 1'h0, _0020_ } | { 1'h0, _0021_ };
  assign _0121_ = - _0263_;
  assign _0123_ = - _0264_;
  assign _0125_ = - _0265_;
  assign _0127_ = - _0266_;
  assign _0122_ = - _0394_;
  assign _0124_ = - _0395_;
  assign _0126_ = - _0396_;
  assign _0128_ = - _0397_;
  assign _0455_ = _0121_ ^ _0122_;
  assign _0456_ = _0123_ ^ _0124_;
  assign _0457_ = _0125_ ^ _0126_;
  assign _0458_ = _0127_ ^ _0128_;
  assign _0502_ = _0455_ | { 27'h0000000, sramreqfifo_rdata_t0[0], 5'h00 };
  assign _0504_ = _0456_ | { 1'h0, _0017_ };
  assign _0506_ = _0457_ | { 1'h0, _0019_ };
  assign _0508_ = _0458_ | { 1'h0, _0021_ };
  assign _0119_ = ~ rspfifo_rvalid;
  assign _0120_ = ~ _0026_;
  assign _0083_ = ~ _0034_;
  assign _0085_ = ~ _0038_;
  assign _0087_ = ~ _0042_;
  assign _0089_ = ~ _0046_;
  assign _0091_ = ~ _0050_;
  assign _0093_ = ~ _0054_;
  assign _0095_ = ~ _0058_;
  assign _0097_ = ~ _0062_;
  assign _0099_ = ~ _0066_;
  assign _0101_ = ~ _0070_;
  assign _0103_ = ~ rspfifo_rdata[0];
  assign _0084_ = ~ { _0032_[23:0], 8'h00 };
  assign _0086_ = ~ { _0036_[23:0], 8'h00 };
  assign _0088_ = ~ { _0040_[15:0], 16'h0000 };
  assign _0090_ = ~ { _0044_[15:0], 16'h0000 };
  assign _0092_ = ~ { _0048_[7:0], 24'h000000 };
  assign _0094_ = ~ { _0052_[7:0], 24'h000000 };
  assign _0096_ = ~ _0000_;
  assign _0098_ = ~ _0002_;
  assign _0100_ = ~ _0004_;
  assign _0102_ = ~ _0006_;
  assign _0267_ = _0035_ & _0084_;
  assign _0270_ = _0039_ & _0086_;
  assign _0273_ = _0043_ & _0088_;
  assign _0276_ = _0047_ & _0090_;
  assign _0279_ = _0051_ & _0092_;
  assign _0282_ = _0055_ & _0094_;
  assign _0285_ = _0059_ & _0096_;
  assign _0288_ = _0063_ & _0098_;
  assign _0291_ = _0067_ & _0100_;
  assign _0294_ = _0071_ & _0102_;
  assign _0297_ = rspfifo_rdata_t0[0] & _0104_;
  assign _0268_ = { _0033_[23:0], 8'h00 } & _0083_;
  assign _0271_ = { _0037_[23:0], 8'h00 } & _0085_;
  assign _0274_ = { _0041_[15:0], 16'h0000 } & _0087_;
  assign _0277_ = { _0045_[15:0], 16'h0000 } & _0089_;
  assign _0280_ = { _0049_[7:0], 24'h000000 } & _0091_;
  assign _0283_ = { _0053_[7:0], 24'h000000 } & _0093_;
  assign _0286_ = _0001_ & _0095_;
  assign _0289_ = _0003_ & _0097_;
  assign _0292_ = _0005_ & _0099_;
  assign _0295_ = _0007_ & _0101_;
  assign _0298_ = reqfifo_rdata_t0[10] & _0103_;
  assign _0269_ = _0035_ & { _0033_[23:0], 8'h00 };
  assign _0272_ = _0039_ & { _0037_[23:0], 8'h00 };
  assign _0275_ = _0043_ & { _0041_[15:0], 16'h0000 };
  assign _0278_ = _0047_ & { _0045_[15:0], 16'h0000 };
  assign _0281_ = _0051_ & { _0049_[7:0], 24'h000000 };
  assign _0284_ = _0055_ & { _0053_[7:0], 24'h000000 };
  assign _0287_ = _0059_ & _0001_;
  assign _0290_ = _0063_ & _0003_;
  assign _0293_ = _0067_ & _0005_;
  assign _0296_ = _0071_ & _0007_;
  assign _0299_ = rspfifo_rdata_t0[0] & reqfifo_rdata_t0[10];
  assign _0398_ = _0267_ | _0268_;
  assign _0399_ = _0270_ | _0271_;
  assign _0400_ = _0273_ | _0274_;
  assign _0401_ = _0276_ | _0277_;
  assign _0402_ = _0279_ | _0280_;
  assign _0403_ = _0282_ | _0283_;
  assign _0404_ = _0285_ | _0286_;
  assign _0405_ = _0288_ | _0289_;
  assign _0406_ = _0291_ | _0292_;
  assign _0407_ = _0294_ | _0295_;
  assign _0408_ = _0297_ | _0298_;
  assign _0515_ = _0398_ | _0269_;
  assign _0517_ = _0399_ | _0272_;
  assign _0519_ = _0400_ | _0275_;
  assign _0521_ = _0401_ | _0278_;
  assign _0522_ = _0402_ | _0281_;
  assign _0523_ = _0403_ | _0284_;
  assign _0525_ = _0404_ | _0287_;
  assign _0527_ = _0405_ | _0290_;
  assign _0529_ = _0406_ | _0293_;
  assign rmask_t0 = _0407_ | _0296_;
  assign _0531_ = _0408_ | _0299_;
  assign _0132_ = | _0502_;
  assign _0133_ = | _0504_;
  assign _0134_ = | _0506_;
  assign _0135_ = | _0508_;
  assign _0471_ = $signed(_0501_) < 0 ? 1'h0 << - _0501_ : 1'h0 >> _0501_;
  assign _0472_ = $signed(_0501_) < 0 ? _0057_ << - _0501_ : _0057_ >> _0501_;
  assign _0473_ = $signed(_0503_) < 0 ? 1'h0 << - _0503_ : 1'h0 >> _0503_;
  assign _0474_ = $signed(_0503_) < 0 ? _0061_ << - _0503_ : _0061_ >> _0503_;
  assign _0475_ = $signed(_0505_) < 0 ? 1'h0 << - _0505_ : 1'h0 >> _0505_;
  assign _0476_ = $signed(_0505_) < 0 ? _0065_ << - _0505_ : _0065_ >> _0505_;
  assign _0477_ = $signed(_0507_) < 0 ? 1'h0 << - _0507_ : 1'h0 >> _0507_;
  assign _0478_ = $signed(_0507_) < 0 ? _0069_ << - _0507_ : _0069_ >> _0507_;
  assign _0009_ = { _0132_, _0132_, _0132_, _0132_, _0132_, _0132_, _0132_, _0132_, _0132_, _0132_, _0132_, _0132_, _0132_, _0132_, _0132_, _0132_, _0132_, _0132_, _0132_, _0132_, _0132_, _0132_, _0132_, _0132_, _0132_, _0132_, _0132_, _0132_, _0132_, _0132_, _0132_, _0132_ } | _0471_;
  assign _0001_ = { _0132_, _0132_, _0132_, _0132_, _0132_, _0132_, _0132_, _0132_, _0132_, _0132_, _0132_, _0132_, _0132_, _0132_, _0132_, _0132_, _0132_, _0132_, _0132_, _0132_, _0132_, _0132_, _0132_, _0132_, _0132_, _0132_, _0132_, _0132_, _0132_, _0132_, _0132_, _0132_ } | _0472_;
  assign _0011_ = { _0133_, _0133_, _0133_, _0133_, _0133_, _0133_, _0133_, _0133_, _0133_, _0133_, _0133_, _0133_, _0133_, _0133_, _0133_, _0133_, _0133_, _0133_, _0133_, _0133_, _0133_, _0133_, _0133_, _0133_, _0133_, _0133_, _0133_, _0133_, _0133_, _0133_, _0133_, _0133_ } | _0473_;
  assign _0003_ = { _0133_, _0133_, _0133_, _0133_, _0133_, _0133_, _0133_, _0133_, _0133_, _0133_, _0133_, _0133_, _0133_, _0133_, _0133_, _0133_, _0133_, _0133_, _0133_, _0133_, _0133_, _0133_, _0133_, _0133_, _0133_, _0133_, _0133_, _0133_, _0133_, _0133_, _0133_, _0133_ } | _0474_;
  assign _0013_ = { _0134_, _0134_, _0134_, _0134_, _0134_, _0134_, _0134_, _0134_, _0134_, _0134_, _0134_, _0134_, _0134_, _0134_, _0134_, _0134_, _0134_, _0134_, _0134_, _0134_, _0134_, _0134_, _0134_, _0134_, _0134_, _0134_, _0134_, _0134_, _0134_, _0134_, _0134_, _0134_ } | _0475_;
  assign _0005_ = { _0134_, _0134_, _0134_, _0134_, _0134_, _0134_, _0134_, _0134_, _0134_, _0134_, _0134_, _0134_, _0134_, _0134_, _0134_, _0134_, _0134_, _0134_, _0134_, _0134_, _0134_, _0134_, _0134_, _0134_, _0134_, _0134_, _0134_, _0134_, _0134_, _0134_, _0134_, _0134_ } | _0476_;
  assign _0015_ = { _0135_, _0135_, _0135_, _0135_, _0135_, _0135_, _0135_, _0135_, _0135_, _0135_, _0135_, _0135_, _0135_, _0135_, _0135_, _0135_, _0135_, _0135_, _0135_, _0135_, _0135_, _0135_, _0135_, _0135_, _0135_, _0135_, _0135_, _0135_, _0135_, _0135_, _0135_, _0135_ } | _0477_;
  assign _0007_ = { _0135_, _0135_, _0135_, _0135_, _0135_, _0135_, _0135_, _0135_, _0135_, _0135_, _0135_, _0135_, _0135_, _0135_, _0135_, _0135_, _0135_, _0135_, _0135_, _0135_, _0135_, _0135_, _0135_, _0135_, _0135_, _0135_, _0135_, _0135_, _0135_, _0135_, _0135_, _0135_ } | _0478_;
  wire [31:0] _1130_ = rdata_t0;
  assign _0479_ = _1130_[$signed({ 26'h0000000, sramreqfifo_rdata[0], 5'h00 }) +: 32];
  assign rdata_tlword_t0 = { sramreqfifo_rdata_t0[0], sramreqfifo_rdata_t0[0], sramreqfifo_rdata_t0[0], sramreqfifo_rdata_t0[0], sramreqfifo_rdata_t0[0], sramreqfifo_rdata_t0[0], sramreqfifo_rdata_t0[0], sramreqfifo_rdata_t0[0], sramreqfifo_rdata_t0[0], sramreqfifo_rdata_t0[0], sramreqfifo_rdata_t0[0], sramreqfifo_rdata_t0[0], sramreqfifo_rdata_t0[0], sramreqfifo_rdata_t0[0], sramreqfifo_rdata_t0[0], sramreqfifo_rdata_t0[0], sramreqfifo_rdata_t0[0], sramreqfifo_rdata_t0[0], sramreqfifo_rdata_t0[0], sramreqfifo_rdata_t0[0], sramreqfifo_rdata_t0[0], sramreqfifo_rdata_t0[0], sramreqfifo_rdata_t0[0], sramreqfifo_rdata_t0[0], sramreqfifo_rdata_t0[0], sramreqfifo_rdata_t0[0], sramreqfifo_rdata_t0[0], sramreqfifo_rdata_t0[0], sramreqfifo_rdata_t0[0], sramreqfifo_rdata_t0[0], sramreqfifo_rdata_t0[0], sramreqfifo_rdata_t0[0] } | _0479_;
  assign _0480_ = reqfifo_rdata[12:11] == 2'h1;
  assign tl_out[1] = d_valid && d_error;
  assign _0482_ = d_valid && _0498_;
  assign _0484_ = d_valid && rspfifo_rvalid;
  assign _0486_ = _0484_ && _0480_;
  assign _0488_ = tl_i[54] && we_o;
  assign _0490_ = tl_i[55] && we_o;
  assign _0492_ = tl_i[56] && we_o;
  assign _0494_ = tl_i[57] && we_o;
  assign _0496_ = ! _0532_;
  assign _0498_ = reqfifo_rdata[12:11] != 2'h1;
  assign _0499_ = tl_i[105:103] != 3'h4;
  assign _0501_ = - $signed({ 27'h0000000, sramreqfifo_rdata[0], 5'h00 });
  assign _0503_ = - $signed({ 1'h0, _0016_ });
  assign _0505_ = - $signed({ 1'h0, _0018_ });
  assign _0507_ = - $signed({ 1'h0, _0020_ });
  assign _0509_ = ~ _0008_;
  assign _0510_ = ~ _0010_;
  assign _0511_ = ~ _0012_;
  assign _0512_ = ~ _0014_;
  assign _0513_ = ~ we_o;
  assign _0514_ = _0034_ | { _0032_[23:0], 8'h00 };
  assign _0516_ = _0038_ | { _0036_[23:0], 8'h00 };
  assign _0518_ = _0042_ | { _0040_[15:0], 16'h0000 };
  assign _0520_ = _0046_ | { _0044_[15:0], 16'h0000 };
  assign _0460_ = _0050_ | { _0048_[7:0], 24'h000000 };
  assign _0459_ = _0054_ | { _0052_[7:0], 24'h000000 };
  assign _0524_ = _0058_ | _0000_;
  assign _0526_ = _0062_ | _0002_;
  assign _0528_ = _0066_ | _0004_;
  assign rmask = _0070_ | _0006_;
  assign _0530_ = rspfifo_rdata[0] | reqfifo_rdata[10];
  assign wdata_o = tl_i[106] ? _0459_ : 32'd0;
  assign wmask_o = tl_i[106] ? _0460_ : 32'd0;
  assign _0022_ = _0480_ ? _0530_ : reqfifo_rdata[10];
  assign d_error = reqfifo_rvalid ? _0022_ : 1'h0;
  assign _0026_ = _0480_ ? rspfifo_rvalid : 1'h1;
  assign _0024_ = reqfifo_rdata[10] ? 1'h1 : _0026_;
  assign d_valid = reqfifo_rvalid ? _0024_ : 1'h0;
  assign _0532_ = | tl_i[105:104];
  assign _0008_ = $signed(_0501_) < 0 ? 8'hff << - _0501_ : 8'hff >> _0501_;
  assign _0000_ = $signed(_0501_) < 0 ? _0056_ << - _0501_ : _0056_ >> _0501_;
  assign _0010_ = $signed(_0503_) < 0 ? 8'hff << - _0503_ : 8'hff >> _0503_;
  assign _0002_ = $signed(_0503_) < 0 ? _0060_ << - _0503_ : _0060_ >> _0503_;
  assign _0012_ = $signed(_0505_) < 0 ? 8'hff << - _0505_ : 8'hff >> _0505_;
  assign _0004_ = $signed(_0505_) < 0 ? _0064_ << - _0505_ : _0064_ >> _0505_;
  assign _0014_ = $signed(_0507_) < 0 ? 8'hff << - _0507_ : 8'hff >> _0507_;
  assign _0006_ = $signed(_0507_) < 0 ? _0068_ << - _0507_ : _0068_ >> _0507_;
  wire [31:0] _1131_ = rdata;
  assign rdata_tlword = _1131_[$signed({ 26'h0000000, sramreqfifo_rdata[0], 5'h00 }) +: 32];
  assign tl_out[64:62] = _0482_ ? 3'h0 : 3'h1;
  assign \sv2v_cast_8DC45$func$generated/sv2v_out.v:9139$90.$result  = d_valid ? rspfifo_rdata[7:1] : 7'h7f;
  assign \sv2v_cast_35AE2$func$generated/sv2v_out.v:9139$93.$result  = _0486_ ? rspfifo_rdata[39:8] : 32'd0;
  assign \sv2v_cast_964CB$func$generated/sv2v_out.v:9139$95.$result  = d_valid ? reqfifo_rdata[7:0] : 8'h00;
  assign \sv2v_cast_4660A$func$generated/sv2v_out.v:9139$96.$result  = d_valid ? reqfifo_rdata[9:8] : 2'h0;
  assign addr_o = tl_i[106] ? tl_i[77:60] : 18'h00000;
  assign _0533_ = _0488_ ? tl_i[29:22] : 8'h00;
  assign _0535_ = _0490_ ? tl_i[37:30] : 8'h00;
  assign _0537_ = _0492_ ? tl_i[45:38] : 8'h00;
  assign _0539_ = _0494_ ? tl_i[53:46] : 8'h00;
  assign reqfifo_wdata[12:11] = _0499_ ? 2'h0 : 2'h1;
  assign rspfifo_rready = _0074_ ? d_ack : 1'h0;
  paramodd4ae9e0467b3ed7a7b38250c0037657e4ca05289auxy_prim_fifo_sync  u_reqfifo (
    .clk_i(clk_i),
    .clr_i(1'h0),
    .clr_i_t0(1'h0),
    .rdata_o(reqfifo_rdata),
    .rdata_o_t0(reqfifo_rdata_t0),
    .rready_i(d_ack),
    .rready_i_t0(d_ack_t0),
    .rst_ni(rst_ni),
    .rvalid_o(reqfifo_rvalid),
    .rvalid_o_t0(reqfifo_rvalid_t0),
    .wdata_i({ reqfifo_wdata[12:11], 1'h0, tl_i[99:90] }),
    .wdata_i_t0({ reqfifo_wdata_t0[12:11], 1'h0, tl_i_t0[99:90] }),
    .wready_o(reqfifo_wready),
    .wready_o_t0(reqfifo_wready_t0),
    .wvalid_i(a_ack),
    .wvalid_i_t0(a_ack_t0)
  );
  paramodauxy_tlul_rsp_intg_genEnableRspIntgGen10EnableDataIntgGen10  u_rsp_gen (
    .tl_i({ d_valid, tl_out[64:62], 3'h0, \sv2v_cast_4660A$func$generated/sv2v_out.v:9139$96.$result , \sv2v_cast_964CB$func$generated/sv2v_out.v:9139$95.$result , 1'h0, \sv2v_cast_35AE2$func$generated/sv2v_out.v:9139$93.$result , 7'h7f, \sv2v_cast_8DC45$func$generated/sv2v_out.v:9139$90.$result , tl_out[1:0] }),
    .tl_i_t0({ d_valid_t0, tl_out_t0[64:62], 3'h0, \sv2v_cast_4660A$func$generated/sv2v_out.v:9139$96.$result_t0 , \sv2v_cast_964CB$func$generated/sv2v_out.v:9139$95.$result_t0 , 1'h0, \sv2v_cast_35AE2$func$generated/sv2v_out.v:9139$93.$result_t0 , 7'h00, \sv2v_cast_8DC45$func$generated/sv2v_out.v:9139$90.$result_t0 , tl_out_t0[1:0] }),
    .tl_o(tl_o),
    .tl_o_t0(tl_o_t0)
  );
  paramoda05994007059a055454376e4d0aa9b8192775615auxy_prim_fifo_sync  u_rspfifo (
    .clk_i(clk_i),
    .clr_i(1'h0),
    .clr_i_t0(1'h0),
    .rdata_o(rspfifo_rdata),
    .rdata_o_t0(rspfifo_rdata_t0),
    .rready_i(rspfifo_rready),
    .rready_i_t0(rspfifo_rready_t0),
    .rst_ni(rst_ni),
    .rvalid_o(rspfifo_rvalid),
    .rvalid_o_t0(rspfifo_rvalid_t0),
    .wdata_i({ rdata_tlword, 7'h7f, rerror_i[1] }),
    .wdata_i_t0({ rdata_tlword_t0, 7'h00, rerror_i_t0[1] }),
    .wready_o(rspfifo_wready),
    .wready_o_t0(rspfifo_wready_t0),
    .wvalid_i(rspfifo_wvalid),
    .wvalid_i_t0(rspfifo_wvalid_t0)
  );
  paramod877a50dace05ef79dab022285c3f67914151b286auxy_prim_fifo_sync  u_sramreqfifo (
    .clk_i(clk_i),
    .clr_i(1'h0),
    .clr_i_t0(1'h0),
    .rdata_o(sramreqfifo_rdata),
    .rdata_o_t0(sramreqfifo_rdata_t0),
    .rready_i(rspfifo_wvalid),
    .rready_i_t0(rspfifo_wvalid_t0),
    .rst_ni(rst_ni),
    .wdata_i({ tl_i[57:54], 1'h0 }),
    .wdata_i_t0({ tl_i_t0[57:54], 1'h0 }),
    .wready_o(sramreqfifo_wready),
    .wready_o_t0(sramreqfifo_wready_t0),
    .wvalid_i(sramreqfifo_wvalid),
    .wvalid_i_t0(sramreqfifo_wvalid_t0)
  );
  assign intg_error_o = 1'h0;
  assign intg_error_o_t0 = 1'h0;
  assign req_type_o = tl_i[16:15];
  assign req_type_o_t0 = tl_i_t0[16:15];
  assign reqfifo_wdata[10:0] = { 1'h0, tl_i[99:90] };
  assign reqfifo_wdata_t0[10:0] = { 1'h0, tl_i_t0[99:90] };
  assign { tl_out[65], tl_out[61:2] } = { d_valid, 3'h0, \sv2v_cast_4660A$func$generated/sv2v_out.v:9139$96.$result , \sv2v_cast_964CB$func$generated/sv2v_out.v:9139$95.$result , 1'h0, \sv2v_cast_35AE2$func$generated/sv2v_out.v:9139$93.$result , 7'h7f, \sv2v_cast_8DC45$func$generated/sv2v_out.v:9139$90.$result  };
  assign { tl_out_t0[65], tl_out_t0[61:2] } = { d_valid_t0, 3'h0, \sv2v_cast_4660A$func$generated/sv2v_out.v:9139$96.$result_t0 , \sv2v_cast_964CB$func$generated/sv2v_out.v:9139$95.$result_t0 , 1'h0, \sv2v_cast_35AE2$func$generated/sv2v_out.v:9139$93.$result_t0 , 7'h00, \sv2v_cast_8DC45$func$generated/sv2v_out.v:9139$90.$result_t0  };
endmodule

module paramodb54d077777a5e0334d1158f40d3ef149c7b94eb9auxy_tlul_fifo_sync (clk_i, rst_ni, tl_h_i, tl_h_o, tl_d_o, tl_d_i, spare_req_i, spare_req_o, spare_rsp_i, spare_rsp_o, spare_rsp_i_t0, spare_req_i_t0, spare_rsp_o_t0, tl_d_i_t0, tl_d_o_t0, tl_h_i_t0, tl_h_o_t0, spare_req_o_t0);
  wire [2:0] _00_;
  wire [31:0] _01_;
  wire _02_;
  wire [2:0] _03_;
  wire [2:0] _04_;
  wire [31:0] _05_;
  wire [31:0] _06_;
  wire [31:0] _07_;
  wire [31:0] _08_;
  wire [31:0] _09_;
  wire [31:0] _10_;
  wire _11_;
  wire _12_;
  wire _13_;
  wire [31:0] _14_;
  wire [31:0] _15_;
  input clk_i;
  wire clk_i;
  input rst_ni;
  wire rst_ni;
  input spare_req_i;
  wire spare_req_i;
  input spare_req_i_t0;
  wire spare_req_i_t0;
  output spare_req_o;
  wire spare_req_o;
  output spare_req_o_t0;
  wire spare_req_o_t0;
  input spare_rsp_i;
  wire spare_rsp_i;
  input spare_rsp_i_t0;
  wire spare_rsp_i_t0;
  output spare_rsp_o;
  wire spare_rsp_o;
  output spare_rsp_o_t0;
  wire spare_rsp_o_t0;
  input [65:0] tl_d_i;
  wire [65:0] tl_d_i;
  input [65:0] tl_d_i_t0;
  wire [65:0] tl_d_i_t0;
  output [106:0] tl_d_o;
  wire [106:0] tl_d_o;
  output [106:0] tl_d_o_t0;
  wire [106:0] tl_d_o_t0;
  input [106:0] tl_h_i;
  wire [106:0] tl_h_i;
  input [106:0] tl_h_i_t0;
  wire [106:0] tl_h_i_t0;
  output [65:0] tl_h_o;
  wire [65:0] tl_h_o;
  output [65:0] tl_h_o_t0;
  wire [65:0] tl_h_o_t0;
  assign _02_ = | tl_d_i_t0[64:62];
  assign _00_ = ~ tl_d_i_t0[64:62];
  assign _03_ = tl_d_i[64:62] & _00_;
  assign _04_ = 3'h1 & _00_;
  assign _11_ = _03_ == _04_;
  assign _13_ = _11_ & _02_;
  assign _01_ = ~ { _12_, _12_, _12_, _12_, _12_, _12_, _12_, _12_, _12_, _12_, _12_, _12_, _12_, _12_, _12_, _12_, _12_, _12_, _12_, _12_, _12_, _12_, _12_, _12_, _12_, _12_, _12_, _12_, _12_, _12_, _12_, _12_ };
  assign _08_ = { _13_, _13_, _13_, _13_, _13_, _13_, _13_, _13_, _13_, _13_, _13_, _13_, _13_, _13_, _13_, _13_, _13_, _13_, _13_, _13_, _13_, _13_, _13_, _13_, _13_, _13_, _13_, _13_, _13_, _13_, _13_, _13_ } | _01_;
  assign _09_ = { _13_, _13_, _13_, _13_, _13_, _13_, _13_, _13_, _13_, _13_, _13_, _13_, _13_, _13_, _13_, _13_, _13_, _13_, _13_, _13_, _13_, _13_, _13_, _13_, _13_, _13_, _13_, _13_, _13_, _13_, _13_, _13_ } | { _12_, _12_, _12_, _12_, _12_, _12_, _12_, _12_, _12_, _12_, _12_, _12_, _12_, _12_, _12_, _12_, _12_, _12_, _12_, _12_, _12_, _12_, _12_, _12_, _12_, _12_, _12_, _12_, _12_, _12_, _12_, _12_ };
  assign _05_ = 32'd0 & _08_;
  assign _06_ = tl_d_i_t0[47:16] & _09_;
  assign _10_ = _05_ | _06_;
  assign _07_ = { _13_, _13_, _13_, _13_, _13_, _13_, _13_, _13_, _13_, _13_, _13_, _13_, _13_, _13_, _13_, _13_, _13_, _13_, _13_, _13_, _13_, _13_, _13_, _13_, _13_, _13_, _13_, _13_, _13_, _13_, _13_, _13_ } & tl_d_i[47:16];
  assign _15_ = _07_ | _10_;
  assign _12_ = tl_d_i[64:62] == 3'h1;
  assign _14_ = _12_ ? tl_d_i[47:16] : 32'd0;
  paramodbcb682b92b2d5f38097d835dce3bd6d5bdad7611auxy_prim_fifo_sync  reqfifo (
    .clk_i(clk_i),
    .clr_i(1'h0),
    .clr_i_t0(1'h0),
    .rdata_o({ tl_d_o[105:1], spare_req_o }),
    .rdata_o_t0({ tl_d_o_t0[105:1], spare_req_o_t0 }),
    .rready_i(tl_d_i[0]),
    .rready_i_t0(tl_d_i_t0[0]),
    .rst_ni(rst_ni),
    .rvalid_o(tl_d_o[106]),
    .rvalid_o_t0(tl_d_o_t0[106]),
    .wdata_i({ tl_h_i[105:1], spare_req_i }),
    .wdata_i_t0({ tl_h_i_t0[105:1], spare_req_i_t0 }),
    .wready_o(tl_h_o[0]),
    .wready_o_t0(tl_h_o_t0[0]),
    .wvalid_i(tl_h_i[106]),
    .wvalid_i_t0(tl_h_i_t0[106])
  );
  paramod4033ffde0d007f439ab68268c14c7a2b914b41b4auxy_prim_fifo_sync  rspfifo (
    .clk_i(clk_i),
    .clr_i(1'h0),
    .clr_i_t0(1'h0),
    .rdata_o({ tl_h_o[64:1], spare_rsp_o }),
    .rdata_o_t0({ tl_h_o_t0[64:1], spare_rsp_o_t0 }),
    .rready_i(tl_h_i[0]),
    .rready_i_t0(tl_h_i_t0[0]),
    .rst_ni(rst_ni),
    .rvalid_o(tl_h_o[65]),
    .rvalid_o_t0(tl_h_o_t0[65]),
    .wdata_i({ tl_d_i[64:48], _14_, tl_d_i[15:1], spare_rsp_i }),
    .wdata_i_t0({ tl_d_i_t0[64:48], _15_, tl_d_i_t0[15:1], spare_rsp_i_t0 }),
    .wready_o(tl_d_o[0]),
    .wready_o_t0(tl_d_o_t0[0]),
    .wvalid_i(tl_d_i[65]),
    .wvalid_i_t0(tl_d_i_t0[65])
  );
endmodule

module paramodbc034ef4e1b4bac0b496e4b04aec5350c1a23f8cauxy_ibex_csr (clk_i, rst_ni, wr_data_i, wr_en_i, rd_data_o, rd_error_o, rd_data_o_t0, rd_error_o_t0, wr_data_i_t0, wr_en_i_t0);
  wire _00_;
  wire _01_;
  wire _02_;
  wire _03_;
  wire _04_;
  wire _05_;
  wire _06_;
  wire _07_;
  wire _08_;
  input clk_i;
  wire clk_i;
  output rd_data_o;
  reg rd_data_o;
  output rd_data_o_t0;
  reg rd_data_o_t0;
  output rd_error_o;
  wire rd_error_o;
  output rd_error_o_t0;
  wire rd_error_o_t0;
  input rst_ni;
  wire rst_ni;
  input wr_data_i;
  wire wr_data_i;
  input wr_data_i_t0;
  wire wr_data_i_t0;
  input wr_en_i;
  wire wr_en_i;
  input wr_en_i_t0;
  wire wr_en_i_t0;
  assign _00_ = ~ wr_en_i;
  assign _08_ = wr_data_i ^ rd_data_o;
  assign _04_ = wr_data_i_t0 | rd_data_o_t0;
  assign _05_ = _08_ | _04_;
  assign _01_ = wr_en_i & wr_data_i_t0;
  assign _02_ = _00_ & rd_data_o_t0;
  assign _03_ = _05_ & wr_en_i_t0;
  assign _06_ = _01_ | _02_;
  assign _07_ = _06_ | _03_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) rd_data_o_t0 <= 1'h0;
    else rd_data_o_t0 <= _07_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) rd_data_o <= 1'h0;
    else if (wr_en_i) rd_data_o <= wr_data_i;
  assign rd_error_o = 1'h0;
  assign rd_error_o_t0 = 1'h0;
endmodule

module paramodbcb682b92b2d5f38097d835dce3bd6d5bdad7611auxy_prim_fifo_sync (clk_i, rst_ni, clr_i, wvalid_i, wready_o, wdata_i, rvalid_o, rready_i, rdata_o, full_o, depth_o, rready_i_t0, rvalid_o_t0, wdata_i_t0, wready_o_t0, wvalid_i_t0, clr_i_t0, depth_o_t0, full_o_t0, rdata_o_t0);
  input clk_i;
  wire clk_i;
  input clr_i;
  wire clr_i;
  input clr_i_t0;
  wire clr_i_t0;
  output depth_o;
  wire depth_o;
  output depth_o_t0;
  wire depth_o_t0;
  output full_o;
  wire full_o;
  output full_o_t0;
  wire full_o_t0;
  output [105:0] rdata_o;
  wire [105:0] rdata_o;
  output [105:0] rdata_o_t0;
  wire [105:0] rdata_o_t0;
  input rready_i;
  wire rready_i;
  input rready_i_t0;
  wire rready_i_t0;
  input rst_ni;
  wire rst_ni;
  output rvalid_o;
  wire rvalid_o;
  output rvalid_o_t0;
  wire rvalid_o_t0;
  input [105:0] wdata_i;
  wire [105:0] wdata_i;
  input [105:0] wdata_i_t0;
  wire [105:0] wdata_i_t0;
  output wready_o;
  wire wready_o;
  output wready_o_t0;
  wire wready_o_t0;
  input wvalid_i;
  wire wvalid_i;
  input wvalid_i_t0;
  wire wvalid_i_t0;
  assign depth_o = 1'h0;
  assign depth_o_t0 = 1'h0;
  assign full_o = rready_i;
  assign full_o_t0 = rready_i_t0;
  assign rdata_o = wdata_i;
  assign rdata_o_t0 = wdata_i_t0;
  assign rvalid_o = wvalid_i;
  assign rvalid_o_t0 = wvalid_i_t0;
  assign wready_o = rready_i;
  assign wready_o_t0 = rready_i_t0;
endmodule

module paramodc28f38d36bce0367a978a541cbb5da157ce66eceauxy_ibex_ex_block (clk_i, rst_ni, alu_operator_i, alu_operand_a_i, alu_operand_b_i, alu_instr_first_cycle_i, bt_a_operand_i, bt_b_operand_i, multdiv_operator_i, mult_en_i, div_en_i, mult_sel_i, div_sel_i, multdiv_signed_mode_i, multdiv_operand_a_i, multdiv_operand_b_i, multdiv_ready_id_i, data_ind_timing_i, imd_val_we_o, imd_val_d_o, imd_val_q_i
, alu_adder_result_ex_o, result_ex_o, branch_target_o, branch_decision_o, ex_valid_o, data_ind_timing_i_t0, imd_val_d_o_t0, imd_val_q_i_t0, imd_val_we_o_t0, multdiv_operand_a_i_t0, multdiv_operand_b_i_t0, div_en_i_t0, div_sel_i_t0, mult_en_i_t0, mult_sel_i_t0, multdiv_ready_id_i_t0, alu_adder_result_ex_o_t0, alu_instr_first_cycle_i_t0, alu_operand_a_i_t0, alu_operand_b_i_t0, alu_operator_i_t0
, branch_decision_o_t0, branch_target_o_t0, bt_a_operand_i_t0, bt_b_operand_i_t0, ex_valid_o_t0, multdiv_operator_i_t0, multdiv_signed_mode_i_t0, result_ex_o_t0);
  wire [32:0] _000_;
  wire [32:0] _001_;
  wire _002_;
  wire _003_;
  wire [1:0] _004_;
  wire [33:0] _005_;
  wire [1:0] _006_;
  wire [31:0] _007_;
  wire _008_;
  wire _009_;
  wire _010_;
  wire [32:0] _011_;
  wire [32:0] _012_;
  wire _013_;
  wire _014_;
  wire _015_;
  wire [1:0] _016_;
  wire [33:0] _017_;
  wire [33:0] _018_;
  wire [33:0] _019_;
  wire [33:0] _020_;
  wire [33:0] _021_;
  wire [33:0] _022_;
  wire [1:0] _023_;
  wire [1:0] _024_;
  wire [1:0] _025_;
  wire [31:0] _026_;
  wire [31:0] _027_;
  wire [31:0] _028_;
  wire _029_;
  wire _030_;
  wire _031_;
  wire [32:0] _032_;
  wire [32:0] _033_;
  wire [32:0] _034_;
  wire _035_;
  wire [33:0] _036_;
  wire [33:0] _037_;
  wire [33:0] _038_;
  wire [33:0] _039_;
  wire [1:0] _040_;
  wire [1:0] _041_;
  wire [1:0] _042_;
  wire [31:0] _043_;
  wire [31:0] _044_;
  wire [31:0] _045_;
  wire _046_;
  wire _047_;
  wire _048_;
  wire [32:0] _049_;
  wire [33:0] _050_;
  wire [33:0] _051_;
  wire [1:0] _052_;
  wire [31:0] _053_;
  wire _054_;
  wire [32:0] _055_;
  wire [32:0] _056_;
  wire _057_;
  wire _058_;
  wire _059_;
  output [31:0] alu_adder_result_ex_o;
  wire [31:0] alu_adder_result_ex_o;
  output [31:0] alu_adder_result_ex_o_t0;
  wire [31:0] alu_adder_result_ex_o_t0;
  wire [33:0] alu_adder_result_ext;
  wire [33:0] alu_adder_result_ext_t0;
  wire [63:0] alu_imd_val_d;
  wire [63:0] alu_imd_val_d_t0;
  wire [1:0] alu_imd_val_we;
  wire [1:0] alu_imd_val_we_t0;
  input alu_instr_first_cycle_i;
  wire alu_instr_first_cycle_i;
  input alu_instr_first_cycle_i_t0;
  wire alu_instr_first_cycle_i_t0;
  wire alu_is_equal_result;
  wire alu_is_equal_result_t0;
  input [31:0] alu_operand_a_i;
  wire [31:0] alu_operand_a_i;
  input [31:0] alu_operand_a_i_t0;
  wire [31:0] alu_operand_a_i_t0;
  input [31:0] alu_operand_b_i;
  wire [31:0] alu_operand_b_i;
  input [31:0] alu_operand_b_i_t0;
  wire [31:0] alu_operand_b_i_t0;
  input [5:0] alu_operator_i;
  wire [5:0] alu_operator_i;
  input [5:0] alu_operator_i_t0;
  wire [5:0] alu_operator_i_t0;
  wire [31:0] alu_result;
  wire [31:0] alu_result_t0;
  output branch_decision_o;
  wire branch_decision_o;
  output branch_decision_o_t0;
  wire branch_decision_o_t0;
  output [31:0] branch_target_o;
  wire [31:0] branch_target_o;
  output [31:0] branch_target_o_t0;
  wire [31:0] branch_target_o_t0;
  input [31:0] bt_a_operand_i;
  wire [31:0] bt_a_operand_i;
  input [31:0] bt_a_operand_i_t0;
  wire [31:0] bt_a_operand_i_t0;
  input [31:0] bt_b_operand_i;
  wire [31:0] bt_b_operand_i;
  input [31:0] bt_b_operand_i_t0;
  wire [31:0] bt_b_operand_i_t0;
  input clk_i;
  wire clk_i;
  input data_ind_timing_i;
  wire data_ind_timing_i;
  input data_ind_timing_i_t0;
  wire data_ind_timing_i_t0;
  input div_en_i;
  wire div_en_i;
  input div_en_i_t0;
  wire div_en_i_t0;
  input div_sel_i;
  wire div_sel_i;
  input div_sel_i_t0;
  wire div_sel_i_t0;
  output ex_valid_o;
  wire ex_valid_o;
  output ex_valid_o_t0;
  wire ex_valid_o_t0;
  wire [32:0] \g_branch_target_alu.bt_alu_result ;
  wire [32:0] \g_branch_target_alu.bt_alu_result_t0 ;
  output [67:0] imd_val_d_o;
  wire [67:0] imd_val_d_o;
  output [67:0] imd_val_d_o_t0;
  wire [67:0] imd_val_d_o_t0;
  input [67:0] imd_val_q_i;
  wire [67:0] imd_val_q_i;
  input [67:0] imd_val_q_i_t0;
  wire [67:0] imd_val_q_i_t0;
  output [1:0] imd_val_we_o;
  wire [1:0] imd_val_we_o;
  output [1:0] imd_val_we_o_t0;
  wire [1:0] imd_val_we_o_t0;
  input mult_en_i;
  wire mult_en_i;
  input mult_en_i_t0;
  wire mult_en_i_t0;
  input mult_sel_i;
  wire mult_sel_i;
  input mult_sel_i_t0;
  wire mult_sel_i_t0;
  wire [32:0] multdiv_alu_operand_a;
  wire [32:0] multdiv_alu_operand_a_t0;
  wire [32:0] multdiv_alu_operand_b;
  wire [32:0] multdiv_alu_operand_b_t0;
  wire [67:0] multdiv_imd_val_d;
  wire [67:0] multdiv_imd_val_d_t0;
  wire [1:0] multdiv_imd_val_we;
  wire [1:0] multdiv_imd_val_we_t0;
  input [31:0] multdiv_operand_a_i;
  wire [31:0] multdiv_operand_a_i;
  input [31:0] multdiv_operand_a_i_t0;
  wire [31:0] multdiv_operand_a_i_t0;
  input [31:0] multdiv_operand_b_i;
  wire [31:0] multdiv_operand_b_i;
  input [31:0] multdiv_operand_b_i_t0;
  wire [31:0] multdiv_operand_b_i_t0;
  input [1:0] multdiv_operator_i;
  wire [1:0] multdiv_operator_i;
  input [1:0] multdiv_operator_i_t0;
  wire [1:0] multdiv_operator_i_t0;
  input multdiv_ready_id_i;
  wire multdiv_ready_id_i;
  input multdiv_ready_id_i_t0;
  wire multdiv_ready_id_i_t0;
  wire [31:0] multdiv_result;
  wire [31:0] multdiv_result_t0;
  wire multdiv_sel;
  wire multdiv_sel_t0;
  input [1:0] multdiv_signed_mode_i;
  wire [1:0] multdiv_signed_mode_i;
  input [1:0] multdiv_signed_mode_i_t0;
  wire [1:0] multdiv_signed_mode_i_t0;
  wire multdiv_valid;
  wire multdiv_valid_t0;
  output [31:0] result_ex_o;
  wire [31:0] result_ex_o;
  output [31:0] result_ex_o_t0;
  wire [31:0] result_ex_o_t0;
  input rst_ni;
  wire rst_ni;
  assign \g_branch_target_alu.bt_alu_result  = bt_a_operand_i + bt_b_operand_i;
  assign _000_ = ~ { 1'h0, bt_a_operand_i_t0 };
  assign _001_ = ~ { 1'h0, bt_b_operand_i_t0 };
  assign _011_ = { 1'h0, bt_a_operand_i } & _000_;
  assign _012_ = { 1'h0, bt_b_operand_i } & _001_;
  assign _055_ = _011_ + _012_;
  assign _032_ = { 1'h0, bt_a_operand_i } | { 1'h0, bt_a_operand_i_t0 };
  assign _033_ = { 1'h0, bt_b_operand_i } | { 1'h0, bt_b_operand_i_t0 };
  assign _056_ = _032_ + _033_;
  assign _049_ = _055_ ^ _056_;
  assign _034_ = _049_ | { 1'h0, bt_a_operand_i_t0 };
  assign \g_branch_target_alu.bt_alu_result_t0  = _034_ | { 1'h0, bt_b_operand_i_t0 };
  assign _009_ = | alu_imd_val_we_t0;
  assign _004_ = ~ alu_imd_val_we_t0;
  assign _016_ = alu_imd_val_we & _004_;
  assign _010_ = ! _016_;
  assign _058_ = _010_ & _009_;
  assign _005_ = ~ { multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel };
  assign _006_ = ~ { multdiv_sel, multdiv_sel };
  assign _007_ = ~ { multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel };
  assign _008_ = ~ multdiv_sel;
  assign _036_ = { multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0 } | _005_;
  assign _040_ = { multdiv_sel_t0, multdiv_sel_t0 } | _006_;
  assign _043_ = { multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0 } | _007_;
  assign _046_ = multdiv_sel_t0 | _008_;
  assign _037_ = { multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0 } | { multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel };
  assign _041_ = { multdiv_sel_t0, multdiv_sel_t0 } | { multdiv_sel, multdiv_sel };
  assign _044_ = { multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0 } | { multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel };
  assign _047_ = multdiv_sel_t0 | multdiv_sel;
  assign _017_ = { 2'h0, alu_imd_val_d_t0[63:32] } & _036_;
  assign _020_ = { 2'h0, alu_imd_val_d_t0[31:0] } & _036_;
  assign _023_ = alu_imd_val_we_t0 & _040_;
  assign _026_ = alu_result_t0 & _043_;
  assign _029_ = _058_ & _046_;
  assign _018_ = multdiv_imd_val_d_t0[67:34] & _037_;
  assign _021_ = multdiv_imd_val_d_t0[33:0] & _037_;
  assign _024_ = multdiv_imd_val_we_t0 & _041_;
  assign _027_ = multdiv_result_t0 & _044_;
  assign _030_ = multdiv_valid_t0 & _047_;
  assign _038_ = _017_ | _018_;
  assign _039_ = _020_ | _021_;
  assign _042_ = _023_ | _024_;
  assign _045_ = _026_ | _027_;
  assign _048_ = _029_ | _030_;
  assign _050_ = { 2'h0, alu_imd_val_d[63:32] } ^ multdiv_imd_val_d[67:34];
  assign _051_ = { 2'h0, alu_imd_val_d[31:0] } ^ multdiv_imd_val_d[33:0];
  assign _052_ = alu_imd_val_we ^ multdiv_imd_val_we;
  assign _053_ = alu_result ^ multdiv_result;
  assign _054_ = _057_ ^ multdiv_valid;
  assign _019_ = { multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0 } & _050_;
  assign _022_ = { multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0 } & _051_;
  assign _025_ = { multdiv_sel_t0, multdiv_sel_t0 } & _052_;
  assign _028_ = { multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0 } & _053_;
  assign _031_ = multdiv_sel_t0 & _054_;
  assign imd_val_d_o_t0[67:34] = _019_ | _038_;
  assign imd_val_d_o_t0[33:0] = _022_ | _039_;
  assign imd_val_we_o_t0 = _025_ | _042_;
  assign result_ex_o_t0 = _028_ | _045_;
  assign ex_valid_o_t0 = _031_ | _048_;
  assign _002_ = ~ mult_sel_i;
  assign _003_ = ~ div_sel_i;
  assign _013_ = mult_sel_i_t0 & _003_;
  assign _014_ = div_sel_i_t0 & _002_;
  assign _015_ = mult_sel_i_t0 & div_sel_i_t0;
  assign _035_ = _013_ | _014_;
  assign multdiv_sel_t0 = _035_ | _015_;
  assign _057_ = ~ _059_;
  assign multdiv_sel = mult_sel_i | div_sel_i;
  assign _059_ = | alu_imd_val_we;
  assign imd_val_d_o[67:34] = multdiv_sel ? multdiv_imd_val_d[67:34] : { 2'h0, alu_imd_val_d[63:32] };
  assign imd_val_d_o[33:0] = multdiv_sel ? multdiv_imd_val_d[33:0] : { 2'h0, alu_imd_val_d[31:0] };
  assign imd_val_we_o = multdiv_sel ? multdiv_imd_val_we : alu_imd_val_we;
  assign result_ex_o = multdiv_sel ? multdiv_result : alu_result;
  assign ex_valid_o = multdiv_sel ? multdiv_valid : _057_;
  paramodauxy_ibex_aluRV32Bs3200000000000000000000000000000000  alu_i (
    .adder_result_ext_o(alu_adder_result_ext),
    .adder_result_ext_o_t0(alu_adder_result_ext_t0),
    .adder_result_o(alu_adder_result_ex_o),
    .adder_result_o_t0(alu_adder_result_ex_o_t0),
    .comparison_result_o(branch_decision_o),
    .comparison_result_o_t0(branch_decision_o_t0),
    .imd_val_d_o(alu_imd_val_d),
    .imd_val_d_o_t0(alu_imd_val_d_t0),
    .imd_val_q_i({ imd_val_q_i[65:34], imd_val_q_i[31:0] }),
    .imd_val_q_i_t0({ imd_val_q_i_t0[65:34], imd_val_q_i_t0[31:0] }),
    .imd_val_we_o(alu_imd_val_we),
    .imd_val_we_o_t0(alu_imd_val_we_t0),
    .instr_first_cycle_i(alu_instr_first_cycle_i),
    .instr_first_cycle_i_t0(alu_instr_first_cycle_i_t0),
    .is_equal_result_o(alu_is_equal_result),
    .is_equal_result_o_t0(alu_is_equal_result_t0),
    .multdiv_operand_a_i(multdiv_alu_operand_a),
    .multdiv_operand_a_i_t0(multdiv_alu_operand_a_t0),
    .multdiv_operand_b_i(multdiv_alu_operand_b),
    .multdiv_operand_b_i_t0(multdiv_alu_operand_b_t0),
    .multdiv_sel_i(multdiv_sel),
    .multdiv_sel_i_t0(multdiv_sel_t0),
    .operand_a_i(alu_operand_a_i),
    .operand_a_i_t0(alu_operand_a_i_t0),
    .operand_b_i(alu_operand_b_i),
    .operand_b_i_t0(alu_operand_b_i_t0),
    .operator_i(alu_operator_i),
    .operator_i_t0(alu_operator_i_t0),
    .result_o(alu_result),
    .result_o_t0(alu_result_t0)
  );
  paramodauxy_ibex_multdiv_fastRV32Ms3200000000000000000000000000000011  \genblk3.gen_multdiv_fast.multdiv_i  (
    .alu_adder_ext_i(alu_adder_result_ext),
    .alu_adder_ext_i_t0(alu_adder_result_ext_t0),
    .alu_adder_i(alu_adder_result_ex_o),
    .alu_adder_i_t0(alu_adder_result_ex_o_t0),
    .alu_operand_a_o(multdiv_alu_operand_a),
    .alu_operand_a_o_t0(multdiv_alu_operand_a_t0),
    .alu_operand_b_o(multdiv_alu_operand_b),
    .alu_operand_b_o_t0(multdiv_alu_operand_b_t0),
    .clk_i(clk_i),
    .data_ind_timing_i(data_ind_timing_i),
    .data_ind_timing_i_t0(data_ind_timing_i_t0),
    .div_en_i(div_en_i),
    .div_en_i_t0(div_en_i_t0),
    .div_sel_i(div_sel_i),
    .div_sel_i_t0(div_sel_i_t0),
    .equal_to_zero_i(alu_is_equal_result),
    .equal_to_zero_i_t0(alu_is_equal_result_t0),
    .imd_val_d_o(multdiv_imd_val_d),
    .imd_val_d_o_t0(multdiv_imd_val_d_t0),
    .imd_val_q_i(imd_val_q_i),
    .imd_val_q_i_t0(imd_val_q_i_t0),
    .imd_val_we_o(multdiv_imd_val_we),
    .imd_val_we_o_t0(multdiv_imd_val_we_t0),
    .mult_en_i(mult_en_i),
    .mult_en_i_t0(mult_en_i_t0),
    .mult_sel_i(mult_sel_i),
    .mult_sel_i_t0(mult_sel_i_t0),
    .multdiv_ready_id_i(multdiv_ready_id_i),
    .multdiv_ready_id_i_t0(multdiv_ready_id_i_t0),
    .multdiv_result_o(multdiv_result),
    .multdiv_result_o_t0(multdiv_result_t0),
    .op_a_i(multdiv_operand_a_i),
    .op_a_i_t0(multdiv_operand_a_i_t0),
    .op_b_i(multdiv_operand_b_i),
    .op_b_i_t0(multdiv_operand_b_i_t0),
    .operator_i(multdiv_operator_i),
    .operator_i_t0(multdiv_operator_i_t0),
    .rst_ni(rst_ni),
    .signed_mode_i(multdiv_signed_mode_i),
    .signed_mode_i_t0(multdiv_signed_mode_i_t0),
    .valid_o(multdiv_valid),
    .valid_o_t0(multdiv_valid_t0)
  );
  assign branch_target_o = \g_branch_target_alu.bt_alu_result [31:0];
  assign branch_target_o_t0 = \g_branch_target_alu.bt_alu_result_t0 [31:0];
endmodule

module paramodc573af43932b4a7bfd8b52400e7bf5041b1b0ddcauxy_ibex_top (clk_i, rst_ni, test_en_i, ram_cfg_i, hart_id_i, boot_addr_i, instr_req_o, instr_gnt_i, instr_rvalid_i, instr_addr_o, instr_rdata_i, instr_err_i, data_req_o, data_gnt_i, data_rvalid_i, data_we_o, data_be_o, data_addr_o, data_wdata_o, data_rdata_i, data_err_i
, irq_software_i, irq_timer_i, irq_external_i, irq_fast_i, irq_nm_i, debug_req_i, crash_dump_o, fetch_enable_i, alert_minor_o, alert_major_o, core_sleep_o, boot_addr_i_t0, test_en_i_t0, instr_rvalid_i_t0, instr_req_o_t0, instr_rdata_i_t0, instr_gnt_i_t0, instr_err_i_t0, instr_addr_o_t0, data_req_o_t0, data_we_o_t0
, debug_req_i_t0, irq_nm_i_t0, data_addr_o_t0, data_be_o_t0, data_err_i_t0, data_gnt_i_t0, data_rdata_i_t0, data_rvalid_i_t0, data_wdata_o_t0, hart_id_i_t0, irq_external_i_t0, irq_fast_i_t0, irq_software_i_t0, irq_timer_i_t0, alert_major_o_t0, alert_minor_o_t0, crash_dump_o_t0, core_sleep_o_t0, fetch_enable_i_t0, ram_cfg_i_t0);
  wire _00_;
  wire _01_;
  wire _02_;
  wire _03_;
  wire _04_;
  wire _05_;
  wire _06_;
  wire _07_;
  wire _08_;
  wire _09_;
  wire _10_;
  wire _11_;
  wire _12_;
  wire _13_;
  wire _14_;
  wire _15_;
  wire _16_;
  wire _17_;
  wire _18_;
  wire _19_;
  wire _20_;
  wire _21_;
  wire _22_;
  wire _23_;
  wire _24_;
  wire _25_;
  wire _26_;
  wire _27_;
  wire _28_;
  wire _29_;
  wire _30_;
  wire _31_;
  wire _32_;
  wire _33_;
  output alert_major_o;
  wire alert_major_o;
  output alert_major_o_t0;
  wire alert_major_o_t0;
  output alert_minor_o;
  wire alert_minor_o;
  output alert_minor_o_t0;
  wire alert_minor_o_t0;
  input [31:0] boot_addr_i;
  wire [31:0] boot_addr_i;
  input [31:0] boot_addr_i_t0;
  wire [31:0] boot_addr_i_t0;
  wire clk;
  input clk_i;
  wire clk_i;
  wire clk_t0;
  wire clock_en;
  wire core_busy_d;
  wire core_busy_d_t0;
  reg core_busy_q;
  reg core_busy_q_t0;
  output core_sleep_o;
  wire core_sleep_o;
  output core_sleep_o_t0;
  wire core_sleep_o_t0;
  output [127:0] crash_dump_o;
  wire [127:0] crash_dump_o;
  output [127:0] crash_dump_o_t0;
  wire [127:0] crash_dump_o_t0;
  output [31:0] data_addr_o;
  wire [31:0] data_addr_o;
  output [31:0] data_addr_o_t0;
  wire [31:0] data_addr_o_t0;
  output [3:0] data_be_o;
  wire [3:0] data_be_o;
  output [3:0] data_be_o_t0;
  wire [3:0] data_be_o_t0;
  input data_err_i;
  wire data_err_i;
  input data_err_i_t0;
  wire data_err_i_t0;
  input data_gnt_i;
  wire data_gnt_i;
  input data_gnt_i_t0;
  wire data_gnt_i_t0;
  input [31:0] data_rdata_i;
  wire [31:0] data_rdata_i;
  input [31:0] data_rdata_i_t0;
  wire [31:0] data_rdata_i_t0;
  output data_req_o;
  wire data_req_o;
  output data_req_o_t0;
  wire data_req_o_t0;
  input data_rvalid_i;
  wire data_rvalid_i;
  input data_rvalid_i_t0;
  wire data_rvalid_i_t0;
  output [31:0] data_wdata_o;
  wire [31:0] data_wdata_o;
  output [31:0] data_wdata_o_t0;
  wire [31:0] data_wdata_o_t0;
  output data_we_o;
  wire data_we_o;
  output data_we_o_t0;
  wire data_we_o_t0;
  input debug_req_i;
  wire debug_req_i;
  input debug_req_i_t0;
  wire debug_req_i_t0;
  wire dummy_instr_id;
  wire dummy_instr_id_t0;
  input fetch_enable_i;
  wire fetch_enable_i;
  input fetch_enable_i_t0;
  wire fetch_enable_i_t0;
  reg fetch_enable_q;
  reg fetch_enable_q_t0;
  input [31:0] hart_id_i;
  wire [31:0] hart_id_i;
  input [31:0] hart_id_i_t0;
  wire [31:0] hart_id_i_t0;
  wire [7:0] ic_data_addr;
  wire [7:0] ic_data_addr_t0;
  wire [1:0] ic_data_req;
  wire [1:0] ic_data_req_t0;
  wire [63:0] ic_data_wdata;
  wire [63:0] ic_data_wdata_t0;
  wire ic_data_write;
  wire ic_data_write_t0;
  wire [7:0] ic_tag_addr;
  wire [7:0] ic_tag_addr_t0;
  wire [1:0] ic_tag_req;
  wire [1:0] ic_tag_req_t0;
  wire [21:0] ic_tag_wdata;
  wire [21:0] ic_tag_wdata_t0;
  wire ic_tag_write;
  wire ic_tag_write_t0;
  output [31:0] instr_addr_o;
  wire [31:0] instr_addr_o;
  output [31:0] instr_addr_o_t0;
  wire [31:0] instr_addr_o_t0;
  input instr_err_i;
  wire instr_err_i;
  input instr_err_i_t0;
  wire instr_err_i_t0;
  input instr_gnt_i;
  wire instr_gnt_i;
  input instr_gnt_i_t0;
  wire instr_gnt_i_t0;
  input [31:0] instr_rdata_i;
  wire [31:0] instr_rdata_i;
  input [31:0] instr_rdata_i_t0;
  wire [31:0] instr_rdata_i_t0;
  output instr_req_o;
  wire instr_req_o;
  output instr_req_o_t0;
  wire instr_req_o_t0;
  input instr_rvalid_i;
  wire instr_rvalid_i;
  input instr_rvalid_i_t0;
  wire instr_rvalid_i_t0;
  input irq_external_i;
  wire irq_external_i;
  input irq_external_i_t0;
  wire irq_external_i_t0;
  input [14:0] irq_fast_i;
  wire [14:0] irq_fast_i;
  input [14:0] irq_fast_i_t0;
  wire [14:0] irq_fast_i_t0;
  input irq_nm_i;
  wire irq_nm_i;
  input irq_nm_i_t0;
  wire irq_nm_i_t0;
  wire irq_pending;
  wire irq_pending_t0;
  input irq_software_i;
  wire irq_software_i;
  input irq_software_i_t0;
  wire irq_software_i_t0;
  input irq_timer_i;
  wire irq_timer_i;
  input irq_timer_i_t0;
  wire irq_timer_i_t0;
  input [9:0] ram_cfg_i;
  wire [9:0] ram_cfg_i;
  input [9:0] ram_cfg_i_t0;
  wire [9:0] ram_cfg_i_t0;
  wire [4:0] rf_raddr_a;
  wire [4:0] rf_raddr_a_t0;
  wire [4:0] rf_raddr_b;
  wire [4:0] rf_raddr_b_t0;
  wire [31:0] rf_rdata_a_ecc;
  wire [31:0] rf_rdata_a_ecc_t0;
  wire [31:0] rf_rdata_b_ecc;
  wire [31:0] rf_rdata_b_ecc_t0;
  wire [4:0] rf_waddr_wb;
  wire [4:0] rf_waddr_wb_t0;
  wire [31:0] rf_wdata_wb_ecc;
  wire [31:0] rf_wdata_wb_ecc_t0;
  wire rf_we_wb;
  wire rf_we_wb_t0;
  input rst_ni;
  wire rst_ni;
  input test_en_i;
  wire test_en_i;
  input test_en_i_t0;
  wire test_en_i_t0;
  assign clock_en = fetch_enable_q & _32_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) core_busy_q_t0 <= 1'h0;
    else core_busy_q_t0 <= core_busy_d_t0;
  assign _00_ = ~ fetch_enable_i;
  assign _23_ = _07_ | fetch_enable_q_t0;
  assign _11_ = _00_ & fetch_enable_q_t0;
  assign _12_ = _23_ & fetch_enable_i_t0;
  assign _24_ = _11_ | _12_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) fetch_enable_q_t0 <= 1'h0;
    else fetch_enable_q_t0 <= _24_;
  assign _08_ = fetch_enable_q_t0 & _32_;
  assign _09_ = _33_ & fetch_enable_q;
  assign _10_ = fetch_enable_q_t0 & _33_;
  assign _22_ = _08_ | _09_;
  assign core_sleep_o_t0 = _22_ | _10_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) fetch_enable_q <= 1'h0;
    else if (fetch_enable_i) fetch_enable_q <= 1'h1;
  assign _07_ = ~ fetch_enable_q;
  assign _01_ = ~ core_busy_q;
  assign _03_ = ~ _28_;
  assign _05_ = ~ _30_;
  assign _02_ = ~ debug_req_i;
  assign _04_ = ~ irq_pending;
  assign _06_ = ~ irq_nm_i;
  assign _13_ = core_busy_q_t0 & _02_;
  assign _16_ = _29_ & _04_;
  assign _19_ = _31_ & _06_;
  assign _14_ = debug_req_i_t0 & _01_;
  assign _17_ = irq_pending_t0 & _03_;
  assign _20_ = irq_nm_i_t0 & _05_;
  assign _15_ = core_busy_q_t0 & debug_req_i_t0;
  assign _18_ = _29_ & irq_pending_t0;
  assign _21_ = _31_ & irq_nm_i_t0;
  assign _25_ = _13_ | _14_;
  assign _26_ = _16_ | _17_;
  assign _27_ = _19_ | _20_;
  assign _29_ = _25_ | _15_;
  assign _31_ = _26_ | _18_;
  assign _33_ = _27_ | _21_;
  assign core_sleep_o = ~ clock_en;
  assign _28_ = core_busy_q | debug_req_i;
  assign _30_ = _28_ | irq_pending;
  assign _32_ = _30_ | irq_nm_i;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) core_busy_q <= 1'h0;
    else core_busy_q <= core_busy_d;
  auxy_prim_clock_gating core_clock_gate_i (
    .clk_i(clk_i),
    .clk_o(clk),
    .clk_o_t0(clk_t0),
    .en_i(clock_en),
    .en_i_t0(core_sleep_o_t0),
    .test_en_i(test_en_i),
    .test_en_i_t0(test_en_i_t0)
  );
  paramod16bd66fd1d1dbd7c4dd1efdb08bf1560b5c5007aauxy_ibex_register_file_ff  \gen_regfile_ff.register_file_i  (
    .clk_i(clk),
    .dummy_instr_id_i(dummy_instr_id),
    .dummy_instr_id_i_t0(dummy_instr_id_t0),
    .raddr_a_i(rf_raddr_a),
    .raddr_a_i_t0(rf_raddr_a_t0),
    .raddr_b_i(rf_raddr_b),
    .raddr_b_i_t0(rf_raddr_b_t0),
    .rdata_a_o(rf_rdata_a_ecc),
    .rdata_a_o_t0(rf_rdata_a_ecc_t0),
    .rdata_b_o(rf_rdata_b_ecc),
    .rdata_b_o_t0(rf_rdata_b_ecc_t0),
    .rst_ni(rst_ni),
    .test_en_i(test_en_i),
    .test_en_i_t0(test_en_i_t0),
    .waddr_a_i(rf_waddr_wb),
    .waddr_a_i_t0(rf_waddr_wb_t0),
    .wdata_a_i(rf_wdata_wb_ecc),
    .wdata_a_i_t0(rf_wdata_wb_ecc_t0),
    .we_a_i(rf_we_wb),
    .we_a_i_t0(rf_we_wb_t0)
  );
  paramod00798253a2da2b158adcde19e501253b4257bf48auxy_ibex_core  u_ibex_core (
    .alert_major_o(alert_major_o),
    .alert_major_o_t0(alert_major_o_t0),
    .alert_minor_o(alert_minor_o),
    .alert_minor_o_t0(alert_minor_o_t0),
    .boot_addr_i(boot_addr_i),
    .boot_addr_i_t0(boot_addr_i_t0),
    .clk_i(clk),
    .core_busy_o(core_busy_d),
    .core_busy_o_t0(core_busy_d_t0),
    .crash_dump_o(crash_dump_o),
    .crash_dump_o_t0(crash_dump_o_t0),
    .data_addr_o(data_addr_o),
    .data_addr_o_t0(data_addr_o_t0),
    .data_be_o(data_be_o),
    .data_be_o_t0(data_be_o_t0),
    .data_err_i(data_err_i),
    .data_err_i_t0(data_err_i_t0),
    .data_gnt_i(data_gnt_i),
    .data_gnt_i_t0(data_gnt_i_t0),
    .data_rdata_i(data_rdata_i),
    .data_rdata_i_t0(data_rdata_i_t0),
    .data_req_o(data_req_o),
    .data_req_o_t0(data_req_o_t0),
    .data_rvalid_i(data_rvalid_i),
    .data_rvalid_i_t0(data_rvalid_i_t0),
    .data_wdata_o(data_wdata_o),
    .data_wdata_o_t0(data_wdata_o_t0),
    .data_we_o(data_we_o),
    .data_we_o_t0(data_we_o_t0),
    .debug_req_i(debug_req_i),
    .debug_req_i_t0(debug_req_i_t0),
    .dummy_instr_id_o(dummy_instr_id),
    .dummy_instr_id_o_t0(dummy_instr_id_t0),
    .hart_id_i(hart_id_i),
    .hart_id_i_t0(hart_id_i_t0),
    .ic_data_addr_o(ic_data_addr),
    .ic_data_addr_o_t0(ic_data_addr_t0),
    .ic_data_rdata_i(128'h00000000000000000000000000000000),
    .ic_data_rdata_i_t0(128'h00000000000000000000000000000000),
    .ic_data_req_o(ic_data_req),
    .ic_data_req_o_t0(ic_data_req_t0),
    .ic_data_wdata_o(ic_data_wdata),
    .ic_data_wdata_o_t0(ic_data_wdata_t0),
    .ic_data_write_o(ic_data_write),
    .ic_data_write_o_t0(ic_data_write_t0),
    .ic_tag_addr_o(ic_tag_addr),
    .ic_tag_addr_o_t0(ic_tag_addr_t0),
    .ic_tag_rdata_i(44'h00000000000),
    .ic_tag_rdata_i_t0(44'h00000000000),
    .ic_tag_req_o(ic_tag_req),
    .ic_tag_req_o_t0(ic_tag_req_t0),
    .ic_tag_wdata_o(ic_tag_wdata),
    .ic_tag_wdata_o_t0(ic_tag_wdata_t0),
    .ic_tag_write_o(ic_tag_write),
    .ic_tag_write_o_t0(ic_tag_write_t0),
    .instr_addr_o(instr_addr_o),
    .instr_addr_o_t0(instr_addr_o_t0),
    .instr_err_i(instr_err_i),
    .instr_err_i_t0(instr_err_i_t0),
    .instr_gnt_i(instr_gnt_i),
    .instr_gnt_i_t0(instr_gnt_i_t0),
    .instr_rdata_i(instr_rdata_i),
    .instr_rdata_i_t0(instr_rdata_i_t0),
    .instr_req_o(instr_req_o),
    .instr_req_o_t0(instr_req_o_t0),
    .instr_rvalid_i(instr_rvalid_i),
    .instr_rvalid_i_t0(instr_rvalid_i_t0),
    .irq_external_i(irq_external_i),
    .irq_external_i_t0(irq_external_i_t0),
    .irq_fast_i(irq_fast_i),
    .irq_fast_i_t0(irq_fast_i_t0),
    .irq_nm_i(irq_nm_i),
    .irq_nm_i_t0(irq_nm_i_t0),
    .irq_pending_o(irq_pending),
    .irq_pending_o_t0(irq_pending_t0),
    .irq_software_i(irq_software_i),
    .irq_software_i_t0(irq_software_i_t0),
    .irq_timer_i(irq_timer_i),
    .irq_timer_i_t0(irq_timer_i_t0),
    .rf_raddr_a_o(rf_raddr_a),
    .rf_raddr_a_o_t0(rf_raddr_a_t0),
    .rf_raddr_b_o(rf_raddr_b),
    .rf_raddr_b_o_t0(rf_raddr_b_t0),
    .rf_rdata_a_ecc_i(rf_rdata_a_ecc),
    .rf_rdata_a_ecc_i_t0(rf_rdata_a_ecc_t0),
    .rf_rdata_b_ecc_i(rf_rdata_b_ecc),
    .rf_rdata_b_ecc_i_t0(rf_rdata_b_ecc_t0),
    .rf_waddr_wb_o(rf_waddr_wb),
    .rf_waddr_wb_o_t0(rf_waddr_wb_t0),
    .rf_wdata_wb_ecc_o(rf_wdata_wb_ecc),
    .rf_wdata_wb_ecc_o_t0(rf_wdata_wb_ecc_t0),
    .rf_we_wb_o(rf_we_wb),
    .rf_we_wb_o_t0(rf_we_wb_t0),
    .rst_ni(rst_ni)
  );
endmodule

module paramodd4ae9e0467b3ed7a7b38250c0037657e4ca05289auxy_prim_fifo_sync (clk_i, rst_ni, clr_i, wvalid_i, wready_o, wdata_i, rvalid_o, rready_i, rdata_o, full_o, depth_o, rready_i_t0, rvalid_o_t0, wdata_i_t0, wready_o_t0, wvalid_i_t0, clr_i_t0, depth_o_t0, full_o_t0, rdata_o_t0);
  wire [1:0] _000_;
  wire [1:0] _001_;
  wire [1:0] _002_;
  wire [1:0] _003_;
  wire _004_;
  wire _005_;
  wire _006_;
  wire _007_;
  wire [1:0] _008_;
  wire [1:0] _009_;
  wire [1:0] _010_;
  wire [1:0] _011_;
  wire _012_;
  wire _013_;
  wire _014_;
  wire _015_;
  wire _016_;
  wire _017_;
  wire _018_;
  wire _019_;
  wire _020_;
  wire _021_;
  wire [1:0] _022_;
  wire [1:0] _023_;
  wire _024_;
  wire _025_;
  wire _026_;
  wire [1:0] _027_;
  wire [1:0] _028_;
  wire _029_;
  wire [1:0] _030_;
  wire [1:0] _031_;
  wire [1:0] _032_;
  wire [1:0] _033_;
  wire [1:0] _034_;
  wire [1:0] _035_;
  wire _036_;
  wire _037_;
  wire _038_;
  wire _039_;
  wire [31:0] _040_;
  wire _041_;
  wire _042_;
  wire _043_;
  wire _044_;
  wire _045_;
  wire _046_;
  wire _047_;
  wire _048_;
  wire _049_;
  wire [1:0] _050_;
  wire [1:0] _051_;
  wire _052_;
  wire _053_;
  wire _054_;
  wire _055_;
  wire _056_;
  wire _057_;
  wire _058_;
  wire _059_;
  wire _060_;
  wire _061_;
  wire _062_;
  wire _063_;
  wire _064_;
  wire _065_;
  wire _066_;
  wire _067_;
  wire _068_;
  wire _069_;
  wire [1:0] _070_;
  wire [1:0] _071_;
  wire [1:0] _072_;
  wire [12:0] _073_;
  wire [12:0] _074_;
  wire [12:0] _075_;
  wire [1:0] _076_;
  wire [1:0] _077_;
  wire [1:0] _078_;
  wire [1:0] _079_;
  wire [1:0] _080_;
  wire _081_;
  wire _082_;
  wire [1:0] _083_;
  wire [1:0] _084_;
  wire [1:0] _085_;
  wire [1:0] _086_;
  wire [1:0] _087_;
  wire [1:0] _088_;
  wire [1:0] _089_;
  wire [1:0] _090_;
  wire [1:0] _091_;
  wire [1:0] _092_;
  wire [1:0] _093_;
  wire [1:0] _094_;
  wire [1:0] _095_;
  wire [1:0] _096_;
  wire [1:0] _097_;
  wire [1:0] _098_;
  wire [1:0] _099_;
  wire [1:0] _100_;
  wire [1:0] _101_;
  wire [1:0] _102_;
  wire _103_;
  wire _104_;
  wire _105_;
  wire _106_;
  wire _107_;
  wire _108_;
  wire _109_;
  wire _110_;
  wire [31:0] _111_;
  wire [31:0] _112_;
  wire [31:0] _113_;
  wire _114_;
  wire _115_;
  wire _116_;
  wire [1:0] _117_;
  wire [1:0] _118_;
  wire _119_;
  wire _120_;
  wire _121_;
  wire _122_;
  wire _123_;
  wire _124_;
  wire [1:0] _125_;
  wire [1:0] _126_;
  wire [1:0] _127_;
  wire [1:0] _128_;
  wire [12:0] _129_;
  wire [12:0] _130_;
  wire [12:0] _131_;
  wire [12:0] _132_;
  wire [1:0] _133_;
  wire [1:0] _134_;
  wire [1:0] _135_;
  wire [1:0] _136_;
  wire _137_;
  wire [1:0] _138_;
  wire [1:0] _139_;
  wire [1:0] _140_;
  wire [1:0] _141_;
  wire [1:0] _142_;
  wire [1:0] _143_;
  wire [1:0] _144_;
  wire [1:0] _145_;
  wire [1:0] _146_;
  wire [1:0] _147_;
  wire [1:0] _148_;
  wire [1:0] _149_;
  wire [1:0] _150_;
  wire [1:0] _151_;
  wire [1:0] _152_;
  wire [1:0] _153_;
  wire [1:0] _154_;
  wire _155_;
  wire _156_;
  wire _157_;
  wire _158_;
  wire _159_;
  wire _160_;
  wire _161_;
  wire _162_;
  wire [31:0] _163_;
  wire [31:0] _164_;
  wire [31:0] _165_;
  wire _166_;
  wire [1:0] _167_;
  wire [1:0] _168_;
  wire [1:0] _169_;
  wire [12:0] _170_;
  wire [1:0] _171_;
  wire [1:0] _172_;
  wire [1:0] _173_;
  wire [1:0] _174_;
  wire [1:0] _175_;
  wire [1:0] _176_;
  wire [1:0] _177_;
  wire _178_;
  wire _179_;
  wire _180_;
  wire _181_;
  wire _182_;
  wire _183_;
  wire _184_;
  wire [1:0] _185_;
  wire [1:0] _186_;
  wire [1:0] _187_;
  wire [1:0] _188_;
  wire _189_;
  wire _190_;
  wire _191_;
  wire _192_;
  wire _193_;
  wire _194_;
  wire _195_;
  wire _196_;
  wire _197_;
  wire [1:0] _198_;
  wire [1:0] _199_;
  wire [1:0] _200_;
  wire [1:0] _201_;
  wire _202_;
  wire _203_;
  wire _204_;
  wire _205_;
  wire _206_;
  wire _207_;
  wire [31:0] _208_;
  wire [31:0] _209_;
  wire [1:0] _210_;
  input clk_i;
  wire clk_i;
  input clr_i;
  wire clr_i;
  input clr_i_t0;
  wire clr_i_t0;
  output depth_o;
  wire depth_o;
  output depth_o_t0;
  wire depth_o_t0;
  output full_o;
  wire full_o;
  output full_o_t0;
  wire full_o_t0;
  wire \gen_normal_fifo.empty ;
  wire \gen_normal_fifo.empty_t0 ;
  wire \gen_normal_fifo.fifo_incr_rptr ;
  wire \gen_normal_fifo.fifo_incr_rptr_t0 ;
  wire \gen_normal_fifo.fifo_incr_wptr ;
  wire \gen_normal_fifo.fifo_incr_wptr_t0 ;
  reg [1:0] \gen_normal_fifo.fifo_rptr ;
  reg [1:0] \gen_normal_fifo.fifo_rptr_t0 ;
  reg [1:0] \gen_normal_fifo.fifo_wptr ;
  reg [1:0] \gen_normal_fifo.fifo_wptr_t0 ;
  reg [12:0] \gen_normal_fifo.rdata_int ;
  reg [12:0] \gen_normal_fifo.rdata_int_t0 ;
  reg \gen_normal_fifo.under_rst ;
  reg \gen_normal_fifo.under_rst_t0 ;
  output [12:0] rdata_o;
  wire [12:0] rdata_o;
  output [12:0] rdata_o_t0;
  wire [12:0] rdata_o_t0;
  input rready_i;
  wire rready_i;
  input rready_i_t0;
  wire rready_i_t0;
  input rst_ni;
  wire rst_ni;
  output rvalid_o;
  wire rvalid_o;
  output rvalid_o_t0;
  wire rvalid_o_t0;
  input [12:0] wdata_i;
  wire [12:0] wdata_i;
  input [12:0] wdata_i_t0;
  wire [12:0] wdata_i_t0;
  output wready_o;
  wire wready_o;
  output wready_o_t0;
  wire wready_o_t0;
  input wvalid_i;
  wire wvalid_i;
  input wvalid_i_t0;
  wire wvalid_i_t0;
  assign _006_ = _204_ + \gen_normal_fifo.fifo_wptr [0];
  assign _008_ = \gen_normal_fifo.fifo_wptr  + 2'h1;
  assign _010_ = \gen_normal_fifo.fifo_rptr  + 2'h1;
  assign _012_ = wvalid_i & wready_o;
  assign \gen_normal_fifo.fifo_incr_wptr  = _012_ & _036_;
  assign _014_ = rvalid_o & rready_i;
  assign \gen_normal_fifo.fifo_incr_rptr  = _014_ & _036_;
  assign wready_o = _039_ & _036_;
  assign rvalid_o = _195_ & _036_;
  assign _020_ = ~ _205_;
  assign _022_ = ~ \gen_normal_fifo.fifo_wptr_t0 ;
  assign _023_ = ~ \gen_normal_fifo.fifo_rptr_t0 ;
  assign _048_ = _204_ & _020_;
  assign _050_ = \gen_normal_fifo.fifo_wptr  & _022_;
  assign _051_ = \gen_normal_fifo.fifo_rptr  & _023_;
  assign _183_ = _048_ + _049_;
  assign _185_ = _050_ + 2'h1;
  assign _187_ = _051_ + 2'h1;
  assign _114_ = _204_ | _205_;
  assign _117_ = \gen_normal_fifo.fifo_wptr  | \gen_normal_fifo.fifo_wptr_t0 ;
  assign _118_ = \gen_normal_fifo.fifo_rptr  | \gen_normal_fifo.fifo_rptr_t0 ;
  assign _184_ = _114_ + _115_;
  assign _186_ = _117_ + 2'h1;
  assign _188_ = _118_ + 2'h1;
  assign _166_ = _183_ ^ _184_;
  assign _167_ = _185_ ^ _186_;
  assign _168_ = _187_ ^ _188_;
  assign _116_ = _166_ | _205_;
  assign _009_ = _167_ | \gen_normal_fifo.fifo_wptr_t0 ;
  assign _011_ = _168_ | \gen_normal_fifo.fifo_rptr_t0 ;
  assign _007_ = _116_ | \gen_normal_fifo.fifo_wptr_t0 [0];
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) \gen_normal_fifo.under_rst_t0  <= 1'h0;
    else \gen_normal_fifo.under_rst_t0  <= _005_;
  assign _024_ = ~ _016_;
  assign _026_ = ~ _018_;
  assign _169_ = _002_ ^ \gen_normal_fifo.fifo_wptr ;
  assign _171_ = _000_ ^ \gen_normal_fifo.fifo_rptr ;
  assign _125_ = _003_ | \gen_normal_fifo.fifo_wptr_t0 ;
  assign _133_ = _001_ | \gen_normal_fifo.fifo_rptr_t0 ;
  assign _126_ = _169_ | _125_;
  assign _134_ = _171_ | _133_;
  assign _070_ = { _016_, _016_ } & _003_;
  assign _076_ = { _018_, _018_ } & _001_;
  assign _071_ = { _024_, _024_ } & \gen_normal_fifo.fifo_wptr_t0 ;
  assign _077_ = { _026_, _026_ } & \gen_normal_fifo.fifo_rptr_t0 ;
  assign _072_ = _126_ & { _017_, _017_ };
  assign _078_ = _134_ & { _019_, _019_ };
  assign _127_ = _070_ | _071_;
  assign _135_ = _076_ | _077_;
  assign _128_ = _127_ | _072_;
  assign _136_ = _135_ | _078_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) \gen_normal_fifo.fifo_wptr_t0  <= 2'h0;
    else \gen_normal_fifo.fifo_wptr_t0  <= _128_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) \gen_normal_fifo.fifo_rptr_t0  <= 2'h0;
    else \gen_normal_fifo.fifo_rptr_t0  <= _136_;
  assign _052_ = wvalid_i_t0 & wready_o;
  assign _055_ = _013_ & _036_;
  assign _058_ = rvalid_o_t0 & rready_i;
  assign _061_ = _015_ & _036_;
  assign _064_ = full_o_t0 & _036_;
  assign _067_ = \gen_normal_fifo.empty_t0  & _036_;
  assign _053_ = wready_o_t0 & wvalid_i;
  assign _056_ = \gen_normal_fifo.under_rst_t0  & _012_;
  assign _059_ = rready_i_t0 & rvalid_o;
  assign _062_ = \gen_normal_fifo.under_rst_t0  & _014_;
  assign _065_ = \gen_normal_fifo.under_rst_t0  & _039_;
  assign _068_ = \gen_normal_fifo.under_rst_t0  & _195_;
  assign _054_ = wvalid_i_t0 & wready_o_t0;
  assign _057_ = _013_ & \gen_normal_fifo.under_rst_t0 ;
  assign _060_ = rvalid_o_t0 & rready_i_t0;
  assign _063_ = _015_ & \gen_normal_fifo.under_rst_t0 ;
  assign _066_ = full_o_t0 & \gen_normal_fifo.under_rst_t0 ;
  assign _069_ = \gen_normal_fifo.empty_t0  & \gen_normal_fifo.under_rst_t0 ;
  assign _119_ = _052_ | _053_;
  assign _120_ = _055_ | _056_;
  assign _121_ = _058_ | _059_;
  assign _122_ = _061_ | _062_;
  assign _123_ = _064_ | _065_;
  assign _124_ = _067_ | _068_;
  assign _013_ = _119_ | _054_;
  assign \gen_normal_fifo.fifo_incr_wptr_t0  = _120_ | _057_;
  assign _015_ = _121_ | _060_;
  assign \gen_normal_fifo.fifo_incr_rptr_t0  = _122_ | _063_;
  assign wready_o_t0 = _123_ | _066_;
  assign rvalid_o_t0 = _124_ | _069_;
  assign _170_ = wdata_i ^ \gen_normal_fifo.rdata_int ;
  assign _025_ = ~ \gen_normal_fifo.fifo_incr_wptr ;
  assign _129_ = wdata_i_t0 | \gen_normal_fifo.rdata_int_t0 ;
  assign _130_ = _170_ | _129_;
  assign _073_ = { \gen_normal_fifo.fifo_incr_wptr , \gen_normal_fifo.fifo_incr_wptr , \gen_normal_fifo.fifo_incr_wptr , \gen_normal_fifo.fifo_incr_wptr , \gen_normal_fifo.fifo_incr_wptr , \gen_normal_fifo.fifo_incr_wptr , \gen_normal_fifo.fifo_incr_wptr , \gen_normal_fifo.fifo_incr_wptr , \gen_normal_fifo.fifo_incr_wptr , \gen_normal_fifo.fifo_incr_wptr , \gen_normal_fifo.fifo_incr_wptr , \gen_normal_fifo.fifo_incr_wptr , \gen_normal_fifo.fifo_incr_wptr  } & wdata_i_t0;
  assign _074_ = { _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_ } & \gen_normal_fifo.rdata_int_t0 ;
  assign _075_ = _130_ & \gen_normal_fifo.fifo_incr_wptr_t0 ;
  assign _131_ = _073_ | _074_;
  assign _132_ = _131_ | _075_;
  always_ff @(posedge clk_i)
    \gen_normal_fifo.rdata_int_t0  <= _132_;
  assign _044_ = | { \gen_normal_fifo.fifo_rptr_t0 [1], \gen_normal_fifo.fifo_wptr_t0 [1] };
  assign _045_ = | { \gen_normal_fifo.fifo_rptr_t0 , \gen_normal_fifo.fifo_wptr_t0  };
  assign _137_ = \gen_normal_fifo.fifo_wptr_t0 [1] | \gen_normal_fifo.fifo_rptr_t0 [1];
  assign _138_ = \gen_normal_fifo.fifo_wptr_t0  | \gen_normal_fifo.fifo_rptr_t0 ;
  assign _029_ = ~ _137_;
  assign _030_ = ~ _138_;
  assign _081_ = \gen_normal_fifo.fifo_wptr [1] & _029_;
  assign _083_ = \gen_normal_fifo.fifo_wptr  & _030_;
  assign _082_ = \gen_normal_fifo.fifo_rptr [1] & _029_;
  assign _084_ = _210_ & _030_;
  assign _085_ = \gen_normal_fifo.fifo_rptr  & _030_;
  assign _180_ = _081_ == _082_;
  assign _181_ = _083_ == _084_;
  assign _182_ = _083_ == _085_;
  assign _194_ = _180_ & _044_;
  assign full_o_t0 = _181_ & _045_;
  assign \gen_normal_fifo.empty_t0  = _182_ & _045_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) \gen_normal_fifo.fifo_wptr  <= 2'h0;
    else if (_016_) \gen_normal_fifo.fifo_wptr  <= _002_;
  always_ff @(posedge clk_i)
    if (\gen_normal_fifo.fifo_incr_wptr ) \gen_normal_fifo.rdata_int  <= wdata_i;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) \gen_normal_fifo.fifo_rptr  <= 2'h0;
    else if (_018_) \gen_normal_fifo.fifo_rptr  <= _000_;
  assign _042_ = | { \gen_normal_fifo.fifo_incr_wptr_t0 , clr_i_t0 };
  assign _043_ = | { \gen_normal_fifo.fifo_incr_rptr_t0 , clr_i_t0 };
  assign _027_ = ~ { \gen_normal_fifo.fifo_incr_wptr_t0 , clr_i_t0 };
  assign _028_ = ~ { \gen_normal_fifo.fifo_incr_rptr_t0 , clr_i_t0 };
  assign _079_ = { \gen_normal_fifo.fifo_incr_wptr , clr_i } & _027_;
  assign _080_ = { \gen_normal_fifo.fifo_incr_rptr , clr_i } & _028_;
  assign _046_ = ! _079_;
  assign _047_ = ! _080_;
  assign _017_ = _046_ & _042_;
  assign _019_ = _047_ & _043_;
  assign _031_ = ~ { \gen_normal_fifo.fifo_rptr [0], \gen_normal_fifo.fifo_rptr [0] };
  assign _032_ = ~ { \gen_normal_fifo.fifo_incr_rptr , \gen_normal_fifo.fifo_incr_rptr  };
  assign _034_ = ~ { \gen_normal_fifo.fifo_wptr [0], \gen_normal_fifo.fifo_wptr [0] };
  assign _035_ = ~ { \gen_normal_fifo.fifo_incr_wptr , \gen_normal_fifo.fifo_incr_wptr  };
  assign _033_ = ~ { clr_i, clr_i };
  assign _036_ = ~ \gen_normal_fifo.under_rst ;
  assign _038_ = ~ _193_;
  assign _039_ = ~ full_o;
  assign _040_ = ~ { \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty  };
  assign _139_ = { \gen_normal_fifo.fifo_rptr_t0 [0], \gen_normal_fifo.fifo_rptr_t0 [0] } | _031_;
  assign _142_ = { \gen_normal_fifo.fifo_incr_rptr_t0 , \gen_normal_fifo.fifo_incr_rptr_t0  } | _032_;
  assign _148_ = { \gen_normal_fifo.fifo_wptr_t0 [0], \gen_normal_fifo.fifo_wptr_t0 [0] } | _034_;
  assign _151_ = { \gen_normal_fifo.fifo_incr_wptr_t0 , \gen_normal_fifo.fifo_incr_wptr_t0  } | _035_;
  assign _145_ = { clr_i_t0, clr_i_t0 } | _033_;
  assign _159_ = _194_ | _038_;
  assign _162_ = full_o_t0 | _039_;
  assign _163_ = { \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0  } | _040_;
  assign _140_ = { \gen_normal_fifo.fifo_rptr_t0 [0], \gen_normal_fifo.fifo_rptr_t0 [0] } | { \gen_normal_fifo.fifo_rptr [0], \gen_normal_fifo.fifo_rptr [0] };
  assign _143_ = { \gen_normal_fifo.fifo_incr_rptr_t0 , \gen_normal_fifo.fifo_incr_rptr_t0  } | { \gen_normal_fifo.fifo_incr_rptr , \gen_normal_fifo.fifo_incr_rptr  };
  assign _149_ = { \gen_normal_fifo.fifo_wptr_t0 [0], \gen_normal_fifo.fifo_wptr_t0 [0] } | { \gen_normal_fifo.fifo_wptr [0], \gen_normal_fifo.fifo_wptr [0] };
  assign _152_ = { \gen_normal_fifo.fifo_incr_wptr_t0 , \gen_normal_fifo.fifo_incr_wptr_t0  } | { \gen_normal_fifo.fifo_incr_wptr , \gen_normal_fifo.fifo_incr_wptr  };
  assign _146_ = { clr_i_t0, clr_i_t0 } | { clr_i, clr_i };
  assign _155_ = \gen_normal_fifo.under_rst_t0  | \gen_normal_fifo.under_rst ;
  assign _160_ = _194_ | _193_;
  assign _164_ = { \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0  } | { \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty , \gen_normal_fifo.empty  };
  assign _086_ = { \gen_normal_fifo.fifo_rptr_t0 [1], 1'h0 } & _139_;
  assign _089_ = 2'h0 & _142_;
  assign _092_ = _199_ & _145_;
  assign _095_ = { \gen_normal_fifo.fifo_wptr_t0 [1], 1'h0 } & _148_;
  assign _098_ = 2'h0 & _151_;
  assign _101_ = _201_ & _145_;
  assign _106_ = _007_ & _159_;
  assign _109_ = _207_ & _162_;
  assign _111_ = { 19'h00000, \gen_normal_fifo.rdata_int_t0  } & _163_;
  assign _087_ = _011_ & _140_;
  assign _090_ = _198_ & _143_;
  assign _096_ = _009_ & _149_;
  assign _099_ = _200_ & _152_;
  assign _093_ = 2'h0 & _146_;
  assign _103_ = \gen_normal_fifo.under_rst_t0  & _155_;
  assign _107_ = _203_ & _160_;
  assign _112_ = 32'd0 & _164_;
  assign _141_ = _086_ | _087_;
  assign _144_ = _089_ | _090_;
  assign _147_ = _092_ | _093_;
  assign _150_ = _095_ | _096_;
  assign _153_ = _098_ | _099_;
  assign _154_ = _101_ | _093_;
  assign _161_ = _106_ | _107_;
  assign _165_ = _111_ | _112_;
  assign _172_ = { _197_, 1'h0 } ^ _010_;
  assign _175_ = { _196_, 1'h0 } ^ _008_;
  assign _179_ = _006_ ^ _202_;
  assign _088_ = { \gen_normal_fifo.fifo_rptr_t0 [0], \gen_normal_fifo.fifo_rptr_t0 [0] } & _172_;
  assign _091_ = { \gen_normal_fifo.fifo_incr_rptr_t0 , \gen_normal_fifo.fifo_incr_rptr_t0  } & _173_;
  assign _094_ = { clr_i_t0, clr_i_t0 } & _174_;
  assign _097_ = { \gen_normal_fifo.fifo_wptr_t0 [0], \gen_normal_fifo.fifo_wptr_t0 [0] } & _175_;
  assign _100_ = { \gen_normal_fifo.fifo_incr_wptr_t0 , \gen_normal_fifo.fifo_incr_wptr_t0  } & _176_;
  assign _102_ = { clr_i_t0, clr_i_t0 } & _177_;
  assign _104_ = \gen_normal_fifo.under_rst_t0  & _036_;
  assign _108_ = _194_ & _179_;
  assign _110_ = full_o_t0 & _041_;
  assign _113_ = { \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0 , \gen_normal_fifo.empty_t0  } & { 19'h00000, \gen_normal_fifo.rdata_int  };
  assign _198_ = _088_ | _141_;
  assign _199_ = _091_ | _144_;
  assign _001_ = _094_ | _147_;
  assign _200_ = _097_ | _150_;
  assign _201_ = _100_ | _153_;
  assign _003_ = _102_ | _154_;
  assign _005_ = _104_ | _103_;
  assign _207_ = _108_ | _161_;
  assign depth_o_t0 = _110_ | _109_;
  assign { _209_[31:13], rdata_o_t0 } = _113_ | _165_;
  assign _016_ = | { \gen_normal_fifo.fifo_incr_wptr , clr_i };
  assign _018_ = | { \gen_normal_fifo.fifo_incr_rptr , clr_i };
  assign _041_ = ~ _206_;
  assign _021_ = ~ \gen_normal_fifo.fifo_wptr_t0 [0];
  assign _037_ = ~ \gen_normal_fifo.fifo_rptr_t0 [0];
  assign _049_ = \gen_normal_fifo.fifo_wptr [0] & _021_;
  assign _105_ = \gen_normal_fifo.fifo_rptr [0] & _037_;
  assign _115_ = \gen_normal_fifo.fifo_wptr [0] | \gen_normal_fifo.fifo_wptr_t0 [0];
  assign _156_ = \gen_normal_fifo.fifo_rptr [0] | \gen_normal_fifo.fifo_rptr_t0 [0];
  assign _189_ = _115_ - _105_;
  assign _191_ = 1'h1 - _105_;
  assign _190_ = _049_ - _156_;
  assign _192_ = 1'h1 - _156_;
  assign _178_ = _189_ ^ _190_;
  assign _158_ = _191_ ^ _192_;
  assign _157_ = _178_ | \gen_normal_fifo.fifo_wptr_t0 [0];
  assign _203_ = _157_ | \gen_normal_fifo.fifo_rptr_t0 [0];
  assign _205_ = _158_ | \gen_normal_fifo.fifo_rptr_t0 [0];
  assign _193_ = \gen_normal_fifo.fifo_wptr [1] == \gen_normal_fifo.fifo_rptr [1];
  assign full_o = \gen_normal_fifo.fifo_wptr  == _210_;
  assign \gen_normal_fifo.empty  = \gen_normal_fifo.fifo_wptr  == \gen_normal_fifo.fifo_rptr ;
  assign _195_ = ~ \gen_normal_fifo.empty ;
  assign _196_ = ~ \gen_normal_fifo.fifo_wptr [1];
  assign _197_ = ~ \gen_normal_fifo.fifo_rptr [1];
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) \gen_normal_fifo.under_rst  <= 1'h1;
    else \gen_normal_fifo.under_rst  <= _004_;
  assign _173_ = \gen_normal_fifo.fifo_rptr [0] ? _010_ : { _197_, 1'h0 };
  assign _174_ = \gen_normal_fifo.fifo_incr_rptr  ? _173_ : 2'hx;
  assign _000_ = clr_i ? 2'h0 : _174_;
  assign _176_ = \gen_normal_fifo.fifo_wptr [0] ? _008_ : { _196_, 1'h0 };
  assign _177_ = \gen_normal_fifo.fifo_incr_wptr  ? _176_ : 2'hx;
  assign _002_ = clr_i ? 2'h0 : _177_;
  assign _004_ = \gen_normal_fifo.under_rst  ? _036_ : 1'h0;
  assign _202_ = \gen_normal_fifo.fifo_wptr [0] - \gen_normal_fifo.fifo_rptr [0];
  assign _204_ = 1'h1 - \gen_normal_fifo.fifo_rptr [0];
  assign _206_ = _193_ ? _202_ : _006_;
  assign depth_o = full_o ? 1'h1 : _206_;
  assign { _208_[31:13], rdata_o } = \gen_normal_fifo.empty  ? 32'd0 : { 19'h00000, \gen_normal_fifo.rdata_int  };
  assign _210_ = \gen_normal_fifo.fifo_rptr  ^ 2'h2;
  assign _208_[12:0] = rdata_o;
  assign _209_[12:0] = rdata_o_t0;
endmodule

module paramode55993a14b1fbc43320d549f521b710ed37596c6auxy_ibex_csr (clk_i, rst_ni, wr_data_i, wr_en_i, rd_data_o, rd_error_o, rd_data_o_t0, rd_error_o_t0, wr_data_i_t0, wr_en_i_t0);
  wire _00_;
  wire [17:0] _01_;
  wire [17:0] _02_;
  wire [17:0] _03_;
  wire [17:0] _04_;
  wire [17:0] _05_;
  wire [17:0] _06_;
  wire [17:0] _07_;
  wire [17:0] _08_;
  input clk_i;
  wire clk_i;
  output [17:0] rd_data_o;
  reg [17:0] rd_data_o;
  output [17:0] rd_data_o_t0;
  reg [17:0] rd_data_o_t0;
  output rd_error_o;
  wire rd_error_o;
  output rd_error_o_t0;
  wire rd_error_o_t0;
  input rst_ni;
  wire rst_ni;
  input [17:0] wr_data_i;
  wire [17:0] wr_data_i;
  input [17:0] wr_data_i_t0;
  wire [17:0] wr_data_i_t0;
  input wr_en_i;
  wire wr_en_i;
  input wr_en_i_t0;
  wire wr_en_i_t0;
  assign _00_ = ~ wr_en_i;
  assign _08_ = wr_data_i ^ rd_data_o;
  assign _04_ = wr_data_i_t0 | rd_data_o_t0;
  assign _05_ = _08_ | _04_;
  assign _01_ = { wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i } & wr_data_i_t0;
  assign _02_ = { _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_ } & rd_data_o_t0;
  assign _03_ = _05_ & { wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0 };
  assign _06_ = _01_ | _02_;
  assign _07_ = _06_ | _03_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) rd_data_o_t0 <= 18'h00000;
    else rd_data_o_t0 <= _07_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) rd_data_o <= 18'h00000;
    else if (wr_en_i) rd_data_o <= wr_data_i;
  assign rd_error_o = 1'h0;
  assign rd_error_o_t0 = 1'h0;
endmodule

module paramode8ca0c7d43bf57ed8b25d9c329a7f7eeb115685cauxy_ibex_id_stage (clk_i, rst_ni, ctrl_busy_o, illegal_insn_o, instr_valid_i, instr_rdata_i, instr_rdata_alu_i, instr_rdata_c_i, instr_is_compressed_i, instr_bp_taken_i, instr_req_o, instr_first_cycle_id_o, instr_valid_clear_o, id_in_ready_o, icache_inval_o, branch_decision_i, pc_set_o, pc_set_spec_o, pc_mux_o, nt_branch_mispredict_o, exc_pc_mux_o
, exc_cause_o, illegal_c_insn_i, instr_fetch_err_i, instr_fetch_err_plus2_i, pc_id_i, ex_valid_i, lsu_resp_valid_i, alu_operator_ex_o, alu_operand_a_ex_o, alu_operand_b_ex_o, imd_val_we_ex_i, imd_val_d_ex_i, imd_val_q_ex_o, bt_a_operand_o, bt_b_operand_o, mult_en_ex_o, div_en_ex_o, mult_sel_ex_o, div_sel_ex_o, multdiv_operator_ex_o, multdiv_signed_mode_ex_o
, multdiv_operand_a_ex_o, multdiv_operand_b_ex_o, multdiv_ready_id_o, csr_access_o, csr_op_o, csr_op_en_o, csr_save_if_o, csr_save_id_o, csr_save_wb_o, csr_restore_mret_id_o, csr_restore_dret_id_o, csr_save_cause_o, csr_mtval_o, priv_mode_i, csr_mstatus_tw_i, illegal_csr_insn_i, data_ind_timing_i, lsu_req_o, lsu_we_o, lsu_type_o, lsu_sign_ext_o
, lsu_wdata_o, lsu_req_done_i, lsu_addr_incr_req_i, lsu_addr_last_i, csr_mstatus_mie_i, irq_pending_i, irqs_i, irq_nm_i, nmi_mode_o, lsu_load_err_i, lsu_store_err_i, debug_mode_o, debug_cause_o, debug_csr_save_o, debug_req_i, debug_single_step_i, debug_ebreakm_i, debug_ebreaku_i, trigger_match_i, result_ex_i, csr_rdata_i
, rf_raddr_a_o, rf_rdata_a_i, rf_raddr_b_o, rf_rdata_b_i, rf_ren_a_o, rf_ren_b_o, rf_waddr_id_o, rf_wdata_id_o, rf_we_id_o, rf_rd_a_wb_match_o, rf_rd_b_wb_match_o, rf_waddr_wb_i, rf_wdata_fwd_wb_i, rf_write_wb_i, en_wb_o, instr_type_wb_o, instr_perf_count_id_o, ready_wb_i, outstanding_load_wb_i, outstanding_store_wb_i, perf_jump_o
, perf_branch_o, perf_tbranch_o, perf_dside_wait_o, perf_mul_wait_o, perf_div_wait_o, instr_id_done_o, instr_req_o_t0, instr_rdata_i_t0, csr_access_o_t0, csr_op_o_t0, icache_inval_o_t0, illegal_insn_o_t0, instr_rdata_alu_i_t0, rf_raddr_a_o_t0, rf_ren_a_o_t0, rf_ren_b_o_t0, rf_raddr_b_o_t0, illegal_c_insn_i_t0, csr_mstatus_mie_i_t0, csr_mstatus_tw_i_t0, csr_mtval_o_t0
, csr_restore_dret_id_o_t0, csr_restore_mret_id_o_t0, csr_save_cause_o_t0, csr_save_id_o_t0, csr_save_if_o_t0, csr_save_wb_o_t0, ctrl_busy_o_t0, debug_cause_o_t0, debug_csr_save_o_t0, debug_ebreakm_i_t0, debug_ebreaku_i_t0, debug_mode_o_t0, debug_req_i_t0, debug_single_step_i_t0, exc_cause_o_t0, exc_pc_mux_o_t0, id_in_ready_o_t0, instr_bp_taken_i_t0, instr_fetch_err_i_t0, instr_fetch_err_plus2_i_t0, instr_is_compressed_i_t0
, instr_valid_clear_o_t0, instr_valid_i_t0, irq_nm_i_t0, irq_pending_i_t0, irqs_i_t0, lsu_addr_last_i_t0, nmi_mode_o_t0, nt_branch_mispredict_o_t0, pc_id_i_t0, pc_mux_o_t0, pc_set_o_t0, pc_set_spec_o_t0, perf_jump_o_t0, perf_tbranch_o_t0, priv_mode_i_t0, ready_wb_i_t0, trigger_match_i_t0, alu_operand_a_ex_o_t0, alu_operand_b_ex_o_t0, alu_operator_ex_o_t0, branch_decision_i_t0
, bt_a_operand_o_t0, bt_b_operand_o_t0, csr_op_en_o_t0, csr_rdata_i_t0, data_ind_timing_i_t0, div_en_ex_o_t0, div_sel_ex_o_t0, en_wb_o_t0, ex_valid_i_t0, illegal_csr_insn_i_t0, imd_val_d_ex_i_t0, imd_val_q_ex_o_t0, imd_val_we_ex_i_t0, instr_first_cycle_id_o_t0, instr_id_done_o_t0, instr_perf_count_id_o_t0, instr_rdata_c_i_t0, instr_type_wb_o_t0, lsu_addr_incr_req_i_t0, lsu_load_err_i_t0, lsu_req_done_i_t0
, lsu_req_o_t0, lsu_resp_valid_i_t0, lsu_sign_ext_o_t0, lsu_store_err_i_t0, lsu_type_o_t0, lsu_wdata_o_t0, lsu_we_o_t0, mult_en_ex_o_t0, mult_sel_ex_o_t0, multdiv_operand_a_ex_o_t0, multdiv_operand_b_ex_o_t0, multdiv_operator_ex_o_t0, multdiv_ready_id_o_t0, multdiv_signed_mode_ex_o_t0, outstanding_load_wb_i_t0, outstanding_store_wb_i_t0, perf_branch_o_t0, perf_div_wait_o_t0, perf_dside_wait_o_t0, perf_mul_wait_o_t0, result_ex_i_t0
, rf_rd_a_wb_match_o_t0, rf_rd_b_wb_match_o_t0, rf_rdata_a_i_t0, rf_rdata_b_i_t0, rf_waddr_id_o_t0, rf_waddr_wb_i_t0, rf_wdata_fwd_wb_i_t0, rf_wdata_id_o_t0, rf_we_id_o_t0, rf_write_wb_i_t0);
  wire _0000_;
  wire _0001_;
  wire _0002_;
  wire _0003_;
  wire _0004_;
  wire _0005_;
  wire _0006_;
  wire _0007_;
  wire _0008_;
  wire _0009_;
  wire _0010_;
  wire _0011_;
  wire _0012_;
  wire _0013_;
  wire _0014_;
  wire _0015_;
  wire _0016_;
  wire _0017_;
  wire _0018_;
  wire _0019_;
  wire _0020_;
  wire _0021_;
  wire _0022_;
  wire _0023_;
  wire _0024_;
  wire _0025_;
  wire _0026_;
  wire _0027_;
  wire _0028_;
  wire _0029_;
  wire _0030_;
  wire _0031_;
  wire _0032_;
  wire _0033_;
  wire _0034_;
  wire _0035_;
  wire _0036_;
  wire _0037_;
  wire _0038_;
  wire _0039_;
  wire _0040_;
  wire _0041_;
  wire _0042_;
  wire _0043_;
  wire _0044_;
  wire _0045_;
  wire _0046_;
  wire _0047_;
  wire _0048_;
  wire _0049_;
  wire _0050_;
  wire _0051_;
  wire _0052_;
  wire _0053_;
  wire _0054_;
  wire _0055_;
  wire _0056_;
  wire _0057_;
  wire _0058_;
  wire _0059_;
  wire _0060_;
  wire _0061_;
  wire _0062_;
  wire _0063_;
  wire _0064_;
  wire _0065_;
  wire _0066_;
  wire _0067_;
  wire _0068_;
  wire _0069_;
  wire _0070_;
  wire _0071_;
  wire _0072_;
  wire _0073_;
  wire _0074_;
  wire _0075_;
  wire _0076_;
  wire _0077_;
  wire _0078_;
  wire _0079_;
  wire _0080_;
  wire _0081_;
  wire _0082_;
  wire _0083_;
  wire _0084_;
  wire _0085_;
  wire _0086_;
  wire _0087_;
  wire _0088_;
  wire _0089_;
  wire _0090_;
  wire _0091_;
  wire _0092_;
  wire _0093_;
  wire _0094_;
  wire _0095_;
  wire _0096_;
  wire _0097_;
  wire _0098_;
  wire _0099_;
  wire _0100_;
  wire _0101_;
  wire [31:0] _0102_;
  wire [31:0] _0103_;
  wire [31:0] _0104_;
  wire [31:0] _0105_;
  wire [31:0] _0106_;
  wire [31:0] _0107_;
  wire [31:0] _0108_;
  wire _0109_;
  wire [31:0] _0110_;
  wire [31:0] _0111_;
  wire [31:0] _0112_;
  wire [31:0] _0113_;
  wire [1:0] _0114_;
  wire [11:0] _0115_;
  wire [4:0] _0116_;
  wire [4:0] _0117_;
  wire _0118_;
  wire _0119_;
  wire _0120_;
  wire _0121_;
  wire _0122_;
  wire _0123_;
  wire _0124_;
  wire _0125_;
  wire _0126_;
  wire _0127_;
  wire _0128_;
  wire _0129_;
  wire _0130_;
  wire _0131_;
  wire _0132_;
  wire _0133_;
  wire _0134_;
  wire _0135_;
  wire _0136_;
  wire _0137_;
  wire _0138_;
  wire _0139_;
  wire _0140_;
  wire _0141_;
  wire _0142_;
  wire _0143_;
  wire _0144_;
  wire _0145_;
  wire _0146_;
  wire _0147_;
  wire _0148_;
  wire _0149_;
  wire _0150_;
  wire _0151_;
  wire _0152_;
  wire _0153_;
  wire _0154_;
  wire _0155_;
  wire [2:0] _0156_;
  wire [2:0] _0157_;
  wire [31:0] _0158_;
  wire [1:0] _0159_;
  wire _0160_;
  wire _0161_;
  wire _0162_;
  wire _0163_;
  wire _0164_;
  wire _0165_;
  wire _0166_;
  wire _0167_;
  wire _0168_;
  wire [1:0] _0169_;
  wire [4:0] _0170_;
  wire [4:0] _0171_;
  wire [1:0] _0172_;
  wire _0173_;
  wire [2:0] _0174_;
  wire [31:0] _0175_;
  wire [31:0] _0176_;
  wire [31:0] _0177_;
  wire [31:0] _0178_;
  wire [31:0] _0179_;
  wire [1:0] _0180_;
  wire [1:0] _0181_;
  wire _0182_;
  wire _0183_;
  wire _0184_;
  wire _0185_;
  wire _0186_;
  wire _0187_;
  wire _0188_;
  wire _0189_;
  wire _0190_;
  wire _0191_;
  wire _0192_;
  wire _0193_;
  wire _0194_;
  wire _0195_;
  wire _0196_;
  wire _0197_;
  wire _0198_;
  wire _0199_;
  wire _0200_;
  wire _0201_;
  wire _0202_;
  wire _0203_;
  wire _0204_;
  wire _0205_;
  wire _0206_;
  wire _0207_;
  wire _0208_;
  wire _0209_;
  wire _0210_;
  wire _0211_;
  wire _0212_;
  wire _0213_;
  wire _0214_;
  wire _0215_;
  wire _0216_;
  wire _0217_;
  wire _0218_;
  wire _0219_;
  wire _0220_;
  wire _0221_;
  wire _0222_;
  wire _0223_;
  wire _0224_;
  wire _0225_;
  wire _0226_;
  wire _0227_;
  wire _0228_;
  wire _0229_;
  wire _0230_;
  wire _0231_;
  wire _0232_;
  wire _0233_;
  wire _0234_;
  wire _0235_;
  wire _0236_;
  wire _0237_;
  wire _0238_;
  wire _0239_;
  wire _0240_;
  wire _0241_;
  wire _0242_;
  wire _0243_;
  wire _0244_;
  wire _0245_;
  wire _0246_;
  wire _0247_;
  wire _0248_;
  wire _0249_;
  wire _0250_;
  wire _0251_;
  wire _0252_;
  wire _0253_;
  wire _0254_;
  wire _0255_;
  wire _0256_;
  wire _0257_;
  wire _0258_;
  wire _0259_;
  wire _0260_;
  wire _0261_;
  wire _0262_;
  wire _0263_;
  wire _0264_;
  wire _0265_;
  wire _0266_;
  wire _0267_;
  wire _0268_;
  wire _0269_;
  wire _0270_;
  wire _0271_;
  wire _0272_;
  wire _0273_;
  wire _0274_;
  wire _0275_;
  wire _0276_;
  wire _0277_;
  wire _0278_;
  wire _0279_;
  wire _0280_;
  wire _0281_;
  wire _0282_;
  wire _0283_;
  wire _0284_;
  wire _0285_;
  wire _0286_;
  wire _0287_;
  wire _0288_;
  wire _0289_;
  wire _0290_;
  wire _0291_;
  wire _0292_;
  wire _0293_;
  wire _0294_;
  wire _0295_;
  wire _0296_;
  wire _0297_;
  wire _0298_;
  wire _0299_;
  wire _0300_;
  wire _0301_;
  wire _0302_;
  wire _0303_;
  wire _0304_;
  wire _0305_;
  wire _0306_;
  wire _0307_;
  wire _0308_;
  wire _0309_;
  wire _0310_;
  wire _0311_;
  wire _0312_;
  wire _0313_;
  wire _0314_;
  wire _0315_;
  wire _0316_;
  wire _0317_;
  wire _0318_;
  wire _0319_;
  wire _0320_;
  wire _0321_;
  wire _0322_;
  wire _0323_;
  wire _0324_;
  wire _0325_;
  wire _0326_;
  wire _0327_;
  wire _0328_;
  wire _0329_;
  wire _0330_;
  wire [33:0] _0331_;
  wire [33:0] _0332_;
  wire [33:0] _0333_;
  wire [33:0] _0334_;
  wire [33:0] _0335_;
  wire [33:0] _0336_;
  wire _0337_;
  wire _0338_;
  wire _0339_;
  wire _0340_;
  wire _0341_;
  wire _0342_;
  wire _0343_;
  wire _0344_;
  wire _0345_;
  wire [31:0] _0346_;
  wire [31:0] _0347_;
  wire [31:0] _0348_;
  wire [31:0] _0349_;
  wire [31:0] _0350_;
  wire [31:0] _0351_;
  wire [31:0] _0352_;
  wire [31:0] _0353_;
  wire [31:0] _0354_;
  wire [31:0] _0355_;
  wire [31:0] _0356_;
  wire [31:0] _0357_;
  wire [31:0] _0358_;
  wire [31:0] _0359_;
  wire [31:0] _0360_;
  wire [31:0] _0361_;
  wire [31:0] _0362_;
  wire [31:0] _0363_;
  wire [31:0] _0364_;
  wire [31:0] _0365_;
  wire [31:0] _0366_;
  wire _0367_;
  wire _0368_;
  wire _0369_;
  wire _0370_;
  wire _0371_;
  wire _0372_;
  wire _0373_;
  wire _0374_;
  wire _0375_;
  wire _0376_;
  wire _0377_;
  wire _0378_;
  wire _0379_;
  wire _0380_;
  wire _0381_;
  wire _0382_;
  wire _0383_;
  wire _0384_;
  wire _0385_;
  wire _0386_;
  wire _0387_;
  wire _0388_;
  wire _0389_;
  wire _0390_;
  wire [31:0] _0391_;
  wire [31:0] _0392_;
  wire [31:0] _0393_;
  wire [31:0] _0394_;
  wire [31:0] _0395_;
  wire [31:0] _0396_;
  wire [31:0] _0397_;
  wire [31:0] _0398_;
  wire [31:0] _0399_;
  wire [31:0] _0400_;
  wire [31:0] _0401_;
  wire [31:0] _0402_;
  wire [1:0] _0403_;
  wire [1:0] _0404_;
  wire [1:0] _0405_;
  wire [11:0] _0406_;
  wire [11:0] _0407_;
  wire [11:0] _0408_;
  wire [11:0] _0409_;
  wire [11:0] _0410_;
  wire [11:0] _0411_;
  wire [11:0] _0412_;
  wire [4:0] _0413_;
  wire [4:0] _0414_;
  wire [4:0] _0415_;
  wire [4:0] _0416_;
  wire _0417_;
  wire _0418_;
  wire _0419_;
  wire _0420_;
  wire _0421_;
  wire _0422_;
  wire _0423_;
  wire _0424_;
  wire _0425_;
  wire _0426_;
  wire _0427_;
  wire _0428_;
  wire _0429_;
  wire _0430_;
  wire _0431_;
  wire _0432_;
  wire _0433_;
  wire _0434_;
  wire _0435_;
  wire _0436_;
  wire _0437_;
  wire _0438_;
  wire _0439_;
  wire _0440_;
  wire _0441_;
  wire _0442_;
  wire _0443_;
  wire _0444_;
  wire _0445_;
  wire _0446_;
  wire _0447_;
  wire _0448_;
  wire _0449_;
  wire _0450_;
  wire _0451_;
  wire _0452_;
  wire _0453_;
  wire _0454_;
  wire _0455_;
  wire _0456_;
  wire _0457_;
  wire _0458_;
  wire _0459_;
  wire _0460_;
  wire _0461_;
  wire _0462_;
  wire _0463_;
  wire _0464_;
  wire _0465_;
  wire _0466_;
  wire _0467_;
  wire _0468_;
  wire _0469_;
  wire _0470_;
  wire _0471_;
  wire _0472_;
  wire _0473_;
  wire _0474_;
  wire _0475_;
  wire _0476_;
  wire _0477_;
  wire _0478_;
  wire _0479_;
  wire _0480_;
  wire _0481_;
  wire _0482_;
  wire _0483_;
  wire _0484_;
  wire _0485_;
  wire [2:0] _0486_;
  wire [2:0] _0487_;
  wire [2:0] _0488_;
  wire [2:0] _0489_;
  wire [2:0] _0490_;
  wire [2:0] _0491_;
  wire [2:0] _0492_;
  wire [31:0] _0493_;
  wire [31:0] _0494_;
  wire [31:0] _0495_;
  wire [1:0] _0496_;
  wire _0497_;
  wire _0498_;
  wire _0499_;
  wire _0500_;
  wire _0501_;
  wire _0502_;
  wire _0503_;
  wire _0504_;
  wire _0505_;
  wire _0506_;
  wire _0507_;
  wire _0508_;
  wire _0509_;
  wire _0510_;
  wire _0511_;
  wire _0512_;
  wire _0513_;
  wire _0514_;
  wire _0515_;
  wire _0516_;
  wire _0517_;
  wire _0518_;
  wire _0519_;
  wire _0520_;
  wire _0521_;
  wire _0522_;
  wire _0523_;
  wire _0524_;
  wire _0525_;
  wire _0526_;
  wire _0527_;
  wire _0528_;
  wire _0529_;
  wire _0530_;
  wire _0531_;
  wire _0532_;
  wire _0533_;
  wire _0534_;
  wire _0535_;
  wire _0536_;
  wire _0537_;
  wire _0538_;
  wire _0539_;
  wire _0540_;
  wire _0541_;
  wire _0542_;
  wire _0543_;
  wire _0544_;
  wire _0545_;
  wire _0546_;
  wire _0547_;
  wire _0548_;
  wire _0549_;
  wire _0550_;
  wire _0551_;
  wire _0552_;
  wire _0553_;
  wire _0554_;
  wire _0555_;
  wire _0556_;
  wire _0557_;
  wire _0558_;
  wire _0559_;
  wire _0560_;
  wire _0561_;
  wire _0562_;
  wire _0563_;
  wire _0564_;
  wire _0565_;
  wire _0566_;
  wire _0567_;
  wire _0568_;
  wire _0569_;
  wire _0570_;
  wire _0571_;
  wire _0572_;
  wire _0573_;
  wire _0574_;
  wire _0575_;
  wire _0576_;
  wire _0577_;
  wire _0578_;
  wire _0579_;
  wire _0580_;
  wire _0581_;
  wire _0582_;
  wire _0583_;
  wire _0584_;
  wire _0585_;
  wire _0586_;
  wire _0587_;
  wire _0588_;
  wire _0589_;
  wire _0590_;
  wire _0591_;
  wire _0592_;
  wire [1:0] _0593_;
  wire [1:0] _0594_;
  wire [1:0] _0595_;
  wire [1:0] _0596_;
  wire [4:0] _0597_;
  wire [4:0] _0598_;
  wire [1:0] _0599_;
  wire [1:0] _0600_;
  wire [1:0] _0601_;
  wire _0602_;
  wire _0603_;
  wire [2:0] _0604_;
  wire [2:0] _0605_;
  wire [2:0] _0606_;
  wire [31:0] _0607_;
  wire [31:0] _0608_;
  wire [31:0] _0609_;
  wire [31:0] _0610_;
  wire [31:0] _0611_;
  wire [31:0] _0612_;
  wire [31:0] _0613_;
  wire [31:0] _0614_;
  wire [31:0] _0615_;
  wire _0616_;
  wire _0617_;
  wire _0618_;
  wire _0619_;
  wire _0620_;
  wire _0621_;
  wire _0622_;
  wire _0623_;
  wire _0624_;
  wire [31:0] _0625_;
  wire [31:0] _0626_;
  wire [31:0] _0627_;
  wire [31:0] _0628_;
  wire [31:0] _0629_;
  wire [31:0] _0630_;
  wire [1:0] _0631_;
  wire [1:0] _0632_;
  wire [1:0] _0633_;
  wire [1:0] _0634_;
  wire [1:0] _0635_;
  wire [1:0] _0636_;
  wire _0637_;
  wire _0638_;
  wire _0639_;
  wire _0640_;
  wire _0641_;
  wire _0642_;
  wire _0643_;
  wire _0644_;
  wire _0645_;
  wire _0646_;
  wire _0647_;
  wire _0648_;
  wire _0649_;
  wire _0650_;
  wire _0651_;
  wire _0652_;
  wire _0653_;
  wire _0654_;
  wire _0655_;
  wire _0656_;
  wire _0657_;
  wire _0658_;
  wire _0659_;
  wire _0660_;
  wire _0661_;
  wire _0662_;
  wire _0663_;
  wire _0664_;
  wire _0665_;
  wire _0666_;
  wire _0667_;
  wire _0668_;
  wire _0669_;
  wire _0670_;
  wire _0671_;
  wire _0672_;
  wire _0673_;
  wire _0674_;
  wire _0675_;
  wire _0676_;
  wire _0677_;
  wire _0678_;
  wire _0679_;
  wire _0680_;
  wire _0681_;
  wire _0682_;
  wire _0683_;
  wire _0684_;
  wire _0685_;
  wire _0686_;
  wire _0687_;
  wire _0688_;
  wire _0689_;
  wire [33:0] _0690_;
  wire [33:0] _0691_;
  wire [33:0] _0692_;
  wire [33:0] _0693_;
  wire [33:0] _0694_;
  wire [33:0] _0695_;
  wire [33:0] _0696_;
  wire [33:0] _0697_;
  wire [1:0] _0698_;
  wire _0699_;
  wire _0700_;
  wire _0701_;
  wire [31:0] _0702_;
  wire [31:0] _0703_;
  wire [31:0] _0704_;
  wire [31:0] _0705_;
  wire [31:0] _0706_;
  wire [31:0] _0707_;
  wire [31:0] _0708_;
  wire [31:0] _0709_;
  wire [31:0] _0710_;
  wire [31:0] _0711_;
  wire [31:0] _0712_;
  wire [31:0] _0713_;
  wire [31:0] _0714_;
  wire [31:0] _0715_;
  wire [31:0] _0716_;
  wire [31:0] _0717_;
  wire [31:0] _0718_;
  wire [31:0] _0719_;
  wire [31:0] _0720_;
  wire [31:0] _0721_;
  wire [31:0] _0722_;
  wire _0723_;
  wire _0724_;
  wire _0725_;
  wire _0726_;
  wire _0727_;
  wire _0728_;
  wire [31:0] _0729_;
  wire [31:0] _0730_;
  wire [31:0] _0731_;
  wire [31:0] _0732_;
  wire [31:0] _0733_;
  wire [31:0] _0734_;
  wire [31:0] _0735_;
  wire [31:0] _0736_;
  wire [31:0] _0737_;
  wire [31:0] _0738_;
  wire [31:0] _0739_;
  wire [31:0] _0740_;
  wire [4:0] _0741_;
  wire [4:0] _0742_;
  wire _0743_;
  wire _0744_;
  wire _0745_;
  wire _0746_;
  wire _0747_;
  wire _0748_;
  wire _0749_;
  wire _0750_;
  wire _0751_;
  wire _0752_;
  wire _0753_;
  wire _0754_;
  wire _0755_;
  wire _0756_;
  wire _0757_;
  wire _0758_;
  wire _0759_;
  wire _0760_;
  wire _0761_;
  wire _0762_;
  wire _0763_;
  wire _0764_;
  wire _0765_;
  wire [31:0] _0766_;
  wire [31:0] _0767_;
  wire [31:0] _0768_;
  wire _0769_;
  wire _0770_;
  wire _0771_;
  wire _0772_;
  wire _0773_;
  wire _0774_;
  wire _0775_;
  wire _0776_;
  wire _0777_;
  wire _0778_;
  wire _0779_;
  wire _0780_;
  wire _0781_;
  wire _0782_;
  wire _0783_;
  wire _0784_;
  wire _0785_;
  wire _0786_;
  wire _0787_;
  wire _0788_;
  wire _0789_;
  wire _0790_;
  wire _0791_;
  wire _0792_;
  wire _0793_;
  wire _0794_;
  wire [1:0] _0795_;
  wire [1:0] _0796_;
  wire [1:0] _0797_;
  wire _0798_;
  wire [2:0] _0799_;
  wire [2:0] _0800_;
  wire [2:0] _0801_;
  wire [31:0] _0802_;
  wire [31:0] _0803_;
  wire [31:0] _0804_;
  wire [31:0] _0805_;
  wire [31:0] _0806_;
  wire [31:0] _0807_;
  wire [31:0] _0808_;
  wire [31:0] _0809_;
  wire [31:0] _0810_;
  wire _0811_;
  wire _0812_;
  wire [31:0] _0813_;
  wire [31:0] _0814_;
  wire [31:0] _0815_;
  wire [31:0] _0816_;
  wire [31:0] _0817_;
  wire [31:0] _0818_;
  wire [1:0] _0819_;
  wire [1:0] _0820_;
  wire [1:0] _0821_;
  wire [1:0] _0822_;
  wire [1:0] _0823_;
  wire [1:0] _0824_;
  wire _0825_;
  wire [33:0] _0826_;
  wire [33:0] _0827_;
  wire [31:0] _0828_;
  wire [31:0] _0829_;
  wire [31:0] _0830_;
  wire [31:0] _0831_;
  wire [31:0] _0832_;
  wire [31:0] _0833_;
  wire [31:0] _0834_;
  wire _0835_;
  wire _0836_;
  wire _0837_;
  wire _0838_;
  wire [31:0] _0839_;
  wire [31:0] _0840_;
  wire [31:0] _0841_;
  wire [31:0] _0842_;
  wire [31:0] _0843_;
  wire _0844_;
  wire _0845_;
  wire _0846_;
  wire _0847_;
  wire _0848_;
  wire _0849_;
  wire _0850_;
  wire _0851_;
  wire _0852_;
  wire _0853_;
  wire _0854_;
  wire _0855_;
  wire _0856_;
  wire _0857_;
  wire _0858_;
  wire _0859_;
  wire _0860_;
  wire _0861_;
  wire _0862_;
  wire _0863_;
  wire _0864_;
  wire _0865_;
  wire _0866_;
  wire _0867_;
  wire _0868_;
  wire _0869_;
  wire _0870_;
  wire [1:0] _0871_;
  wire [2:0] _0872_;
  wire [31:0] _0873_;
  wire _0874_;
  wire [31:0] _0875_;
  wire [31:0] _0876_;
  wire [1:0] _0877_;
  wire _0878_;
  wire _0879_;
  wire _0880_;
  wire _0881_;
  wire _0882_;
  wire _0883_;
  wire _0884_;
  wire _0885_;
  wire _0886_;
  wire _0887_;
  wire _0888_;
  wire _0889_;
  wire _0890_;
  wire _0891_;
  wire _0892_;
  wire _0893_;
  wire _0894_;
  wire _0895_;
  wire [31:0] _0896_;
  wire [31:0] _0897_;
  wire [31:0] _0898_;
  wire [31:0] _0899_;
  wire [31:0] _0900_;
  wire [31:0] _0901_;
  wire [31:0] _0902_;
  wire [31:0] _0903_;
  wire [31:0] _0904_;
  wire [31:0] _0905_;
  wire [31:0] _0906_;
  wire [31:0] _0907_;
  wire [31:0] _0908_;
  wire [31:0] _0909_;
  wire _0910_;
  wire _0911_;
  wire _0912_;
  wire _0913_;
  wire _0914_;
  wire _0915_;
  wire _0916_;
  wire _0917_;
  wire _0918_;
  wire _0919_;
  wire _0920_;
  wire _0921_;
  wire _0922_;
  wire _0923_;
  wire _0924_;
  wire _0925_;
  wire _0926_;
  wire _0927_;
  wire _0928_;
  wire _0929_;
  wire _0930_;
  wire _0931_;
  wire _0932_;
  wire _0933_;
  wire _0934_;
  wire _0935_;
  wire _0936_;
  wire _0937_;
  wire _0938_;
  wire _0939_;
  wire _0940_;
  wire _0941_;
  wire _0942_;
  wire _0943_;
  wire _0944_;
  wire _0945_;
  wire _0946_;
  wire _0947_;
  wire _0948_;
  wire _0949_;
  wire _0950_;
  wire _0951_;
  wire _0952_;
  wire _0953_;
  wire _0954_;
  wire _0955_;
  wire _0956_;
  wire _0957_;
  wire _0958_;
  wire _0959_;
  wire _0960_;
  wire _0961_;
  wire _0962_;
  wire _0963_;
  wire _0964_;
  wire _0965_;
  wire _0966_;
  wire _0967_;
  wire _0968_;
  wire _0969_;
  wire _0970_;
  wire _0971_;
  wire _0972_;
  wire _0973_;
  wire _0974_;
  wire _0975_;
  wire _0976_;
  wire _0977_;
  wire _0978_;
  wire _0979_;
  wire _0980_;
  wire _0981_;
  wire _0982_;
  wire _0983_;
  wire _0984_;
  wire _0985_;
  wire _0986_;
  wire _0987_;
  wire _0988_;
  wire _0989_;
  wire _0990_;
  wire _0991_;
  wire _0992_;
  wire _0993_;
  wire _0994_;
  wire _0995_;
  wire _0996_;
  wire _0997_;
  wire _0998_;
  wire _0999_;
  wire _1000_;
  wire _1001_;
  wire _1002_;
  wire _1003_;
  wire _1004_;
  wire _1005_;
  wire _1006_;
  wire _1007_;
  wire _1008_;
  wire _1009_;
  wire _1010_;
  wire _1011_;
  wire _1012_;
  wire _1013_;
  wire _1014_;
  wire _1015_;
  wire _1016_;
  wire _1017_;
  wire _1018_;
  wire _1019_;
  wire _1020_;
  wire _1021_;
  wire _1022_;
  wire _1023_;
  wire _1024_;
  wire _1025_;
  wire _1026_;
  wire _1027_;
  wire _1028_;
  wire _1029_;
  wire _1030_;
  wire [31:0] _1031_;
  wire [31:0] _1032_;
  wire _1033_;
  wire [1:0] _1034_;
  wire [1:0] _1035_;
  wire alu_multicycle_dec;
  wire alu_multicycle_dec_t0;
  wire [1:0] alu_op_a_mux_sel;
  wire [1:0] alu_op_a_mux_sel_dec;
  wire [1:0] alu_op_a_mux_sel_dec_t0;
  wire [1:0] alu_op_a_mux_sel_t0;
  wire alu_op_b_mux_sel;
  wire alu_op_b_mux_sel_dec;
  wire alu_op_b_mux_sel_dec_t0;
  wire alu_op_b_mux_sel_t0;
  output [31:0] alu_operand_a_ex_o;
  wire [31:0] alu_operand_a_ex_o;
  output [31:0] alu_operand_a_ex_o_t0;
  wire [31:0] alu_operand_a_ex_o_t0;
  output [31:0] alu_operand_b_ex_o;
  wire [31:0] alu_operand_b_ex_o;
  output [31:0] alu_operand_b_ex_o_t0;
  wire [31:0] alu_operand_b_ex_o_t0;
  output [5:0] alu_operator_ex_o;
  wire [5:0] alu_operator_ex_o;
  output [5:0] alu_operator_ex_o_t0;
  wire [5:0] alu_operator_ex_o_t0;
  input branch_decision_i;
  wire branch_decision_i;
  input branch_decision_i_t0;
  wire branch_decision_i_t0;
  wire branch_in_dec;
  wire branch_in_dec_t0;
  wire branch_jump_set_done_d;
  wire branch_jump_set_done_d_t0;
  reg branch_jump_set_done_q;
  reg branch_jump_set_done_q_t0;
  wire branch_set;
  wire branch_set_raw;
  wire branch_set_raw_spec;
  wire branch_set_raw_spec_t0;
  wire branch_set_raw_t0;
  wire branch_set_spec;
  wire branch_set_spec_t0;
  wire branch_set_t0;
  wire [1:0] bt_a_mux_sel;
  wire [1:0] bt_a_mux_sel_t0;
  output [31:0] bt_a_operand_o;
  wire [31:0] bt_a_operand_o;
  output [31:0] bt_a_operand_o_t0;
  wire [31:0] bt_a_operand_o_t0;
  wire [2:0] bt_b_mux_sel;
  wire [2:0] bt_b_mux_sel_t0;
  output [31:0] bt_b_operand_o;
  wire [31:0] bt_b_operand_o;
  output [31:0] bt_b_operand_o_t0;
  wire [31:0] bt_b_operand_o_t0;
  input clk_i;
  wire clk_i;
  wire controller_run;
  wire controller_run_t0;
  output csr_access_o;
  wire csr_access_o;
  output csr_access_o_t0;
  wire csr_access_o_t0;
  input csr_mstatus_mie_i;
  wire csr_mstatus_mie_i;
  input csr_mstatus_mie_i_t0;
  wire csr_mstatus_mie_i_t0;
  input csr_mstatus_tw_i;
  wire csr_mstatus_tw_i;
  input csr_mstatus_tw_i_t0;
  wire csr_mstatus_tw_i_t0;
  output [31:0] csr_mtval_o;
  wire [31:0] csr_mtval_o;
  output [31:0] csr_mtval_o_t0;
  wire [31:0] csr_mtval_o_t0;
  output csr_op_en_o;
  wire csr_op_en_o;
  output csr_op_en_o_t0;
  wire csr_op_en_o_t0;
  output [1:0] csr_op_o;
  wire [1:0] csr_op_o;
  output [1:0] csr_op_o_t0;
  wire [1:0] csr_op_o_t0;
  wire csr_pipe_flush;
  wire csr_pipe_flush_t0;
  input [31:0] csr_rdata_i;
  wire [31:0] csr_rdata_i;
  input [31:0] csr_rdata_i_t0;
  wire [31:0] csr_rdata_i_t0;
  output csr_restore_dret_id_o;
  wire csr_restore_dret_id_o;
  output csr_restore_dret_id_o_t0;
  wire csr_restore_dret_id_o_t0;
  output csr_restore_mret_id_o;
  wire csr_restore_mret_id_o;
  output csr_restore_mret_id_o_t0;
  wire csr_restore_mret_id_o_t0;
  output csr_save_cause_o;
  wire csr_save_cause_o;
  output csr_save_cause_o_t0;
  wire csr_save_cause_o_t0;
  output csr_save_id_o;
  wire csr_save_id_o;
  output csr_save_id_o_t0;
  wire csr_save_id_o_t0;
  output csr_save_if_o;
  wire csr_save_if_o;
  output csr_save_if_o_t0;
  wire csr_save_if_o_t0;
  output csr_save_wb_o;
  wire csr_save_wb_o;
  output csr_save_wb_o_t0;
  wire csr_save_wb_o_t0;
  output ctrl_busy_o;
  wire ctrl_busy_o;
  output ctrl_busy_o_t0;
  wire ctrl_busy_o_t0;
  input data_ind_timing_i;
  wire data_ind_timing_i;
  input data_ind_timing_i_t0;
  wire data_ind_timing_i_t0;
  wire data_req_allowed;
  wire data_req_allowed_t0;
  output [2:0] debug_cause_o;
  wire [2:0] debug_cause_o;
  output [2:0] debug_cause_o_t0;
  wire [2:0] debug_cause_o_t0;
  output debug_csr_save_o;
  wire debug_csr_save_o;
  output debug_csr_save_o_t0;
  wire debug_csr_save_o_t0;
  input debug_ebreakm_i;
  wire debug_ebreakm_i;
  input debug_ebreakm_i_t0;
  wire debug_ebreakm_i_t0;
  input debug_ebreaku_i;
  wire debug_ebreaku_i;
  input debug_ebreaku_i_t0;
  wire debug_ebreaku_i_t0;
  output debug_mode_o;
  wire debug_mode_o;
  output debug_mode_o_t0;
  wire debug_mode_o_t0;
  input debug_req_i;
  wire debug_req_i;
  input debug_req_i_t0;
  wire debug_req_i_t0;
  input debug_single_step_i;
  wire debug_single_step_i;
  input debug_single_step_i_t0;
  wire debug_single_step_i_t0;
  wire div_en_dec;
  wire div_en_dec_t0;
  output div_en_ex_o;
  wire div_en_ex_o;
  output div_en_ex_o_t0;
  wire div_en_ex_o_t0;
  output div_sel_ex_o;
  wire div_sel_ex_o;
  output div_sel_ex_o_t0;
  wire div_sel_ex_o_t0;
  wire dret_insn_dec;
  wire dret_insn_dec_t0;
  wire ebrk_insn;
  wire ebrk_insn_t0;
  wire ecall_insn_dec;
  wire ecall_insn_dec_t0;
  output en_wb_o;
  wire en_wb_o;
  output en_wb_o_t0;
  wire en_wb_o_t0;
  input ex_valid_i;
  wire ex_valid_i;
  input ex_valid_i_t0;
  wire ex_valid_i_t0;
  output [5:0] exc_cause_o;
  wire [5:0] exc_cause_o;
  output [5:0] exc_cause_o_t0;
  wire [5:0] exc_cause_o_t0;
  output [1:0] exc_pc_mux_o;
  wire [1:0] exc_pc_mux_o;
  output [1:0] exc_pc_mux_o_t0;
  wire [1:0] exc_pc_mux_o_t0;
  wire flush_id;
  wire flush_id_t0;
  wire \gen_stall_mem.instr_kill ;
  wire \gen_stall_mem.instr_kill_t0 ;
  wire \gen_stall_mem.outstanding_memory_access ;
  wire \gen_stall_mem.rf_rd_a_hz ;
  wire \gen_stall_mem.rf_rd_a_hz_t0 ;
  wire \gen_stall_mem.rf_rd_b_hz ;
  wire \gen_stall_mem.rf_rd_b_hz_t0 ;
  output icache_inval_o;
  wire icache_inval_o;
  output icache_inval_o_t0;
  wire icache_inval_o_t0;
  reg id_fsm_q;
  reg id_fsm_q_t0;
  output id_in_ready_o;
  wire id_in_ready_o;
  output id_in_ready_o_t0;
  wire id_in_ready_o_t0;
  input illegal_c_insn_i;
  wire illegal_c_insn_i;
  input illegal_c_insn_i_t0;
  wire illegal_c_insn_i_t0;
  input illegal_csr_insn_i;
  wire illegal_csr_insn_i;
  input illegal_csr_insn_i_t0;
  wire illegal_csr_insn_i_t0;
  wire illegal_insn_dec;
  wire illegal_insn_dec_t0;
  output illegal_insn_o;
  wire illegal_insn_o;
  output illegal_insn_o_t0;
  wire illegal_insn_o_t0;
  input [67:0] imd_val_d_ex_i;
  wire [67:0] imd_val_d_ex_i;
  input [67:0] imd_val_d_ex_i_t0;
  wire [67:0] imd_val_d_ex_i_t0;
  output [67:0] imd_val_q_ex_o;
  reg [67:0] imd_val_q_ex_o;
  output [67:0] imd_val_q_ex_o_t0;
  reg [67:0] imd_val_q_ex_o_t0;
  input [1:0] imd_val_we_ex_i;
  wire [1:0] imd_val_we_ex_i;
  input [1:0] imd_val_we_ex_i_t0;
  wire [1:0] imd_val_we_ex_i_t0;
  wire [31:0] imm_a;
  wire imm_a_mux_sel;
  wire imm_a_mux_sel_t0;
  wire [31:0] imm_a_t0;
  wire [31:0] imm_b;
  wire [2:0] imm_b_mux_sel;
  wire [2:0] imm_b_mux_sel_dec;
  wire [2:0] imm_b_mux_sel_dec_t0;
  wire [2:0] imm_b_mux_sel_t0;
  wire [31:0] imm_b_t0;
  wire [31:0] imm_b_type;
  wire [31:0] imm_b_type_t0;
  wire [31:0] imm_i_type;
  wire [31:0] imm_i_type_t0;
  wire [31:0] imm_j_type;
  wire [31:0] imm_j_type_t0;
  wire [31:0] imm_s_type;
  wire [31:0] imm_s_type_t0;
  wire [31:0] imm_u_type;
  wire [31:0] imm_u_type_t0;
  input instr_bp_taken_i;
  wire instr_bp_taken_i;
  input instr_bp_taken_i_t0;
  wire instr_bp_taken_i_t0;
  wire instr_executing;
  wire instr_executing_spec;
  wire instr_executing_spec_t0;
  wire instr_executing_t0;
  input instr_fetch_err_i;
  wire instr_fetch_err_i;
  input instr_fetch_err_i_t0;
  wire instr_fetch_err_i_t0;
  input instr_fetch_err_plus2_i;
  wire instr_fetch_err_plus2_i;
  input instr_fetch_err_plus2_i_t0;
  wire instr_fetch_err_plus2_i_t0;
  output instr_first_cycle_id_o;
  wire instr_first_cycle_id_o;
  output instr_first_cycle_id_o_t0;
  wire instr_first_cycle_id_o_t0;
  output instr_id_done_o;
  wire instr_id_done_o;
  output instr_id_done_o_t0;
  wire instr_id_done_o_t0;
  input instr_is_compressed_i;
  wire instr_is_compressed_i;
  input instr_is_compressed_i_t0;
  wire instr_is_compressed_i_t0;
  output instr_perf_count_id_o;
  wire instr_perf_count_id_o;
  output instr_perf_count_id_o_t0;
  wire instr_perf_count_id_o_t0;
  input [31:0] instr_rdata_alu_i;
  wire [31:0] instr_rdata_alu_i;
  input [31:0] instr_rdata_alu_i_t0;
  wire [31:0] instr_rdata_alu_i_t0;
  input [15:0] instr_rdata_c_i;
  wire [15:0] instr_rdata_c_i;
  input [15:0] instr_rdata_c_i_t0;
  wire [15:0] instr_rdata_c_i_t0;
  input [31:0] instr_rdata_i;
  wire [31:0] instr_rdata_i;
  input [31:0] instr_rdata_i_t0;
  wire [31:0] instr_rdata_i_t0;
  output instr_req_o;
  wire instr_req_o;
  output instr_req_o_t0;
  wire instr_req_o_t0;
  output [1:0] instr_type_wb_o;
  wire [1:0] instr_type_wb_o;
  output [1:0] instr_type_wb_o_t0;
  wire [1:0] instr_type_wb_o_t0;
  output instr_valid_clear_o;
  wire instr_valid_clear_o;
  output instr_valid_clear_o_t0;
  wire instr_valid_clear_o_t0;
  input instr_valid_i;
  wire instr_valid_i;
  input instr_valid_i_t0;
  wire instr_valid_i_t0;
  input irq_nm_i;
  wire irq_nm_i;
  input irq_nm_i_t0;
  wire irq_nm_i_t0;
  input irq_pending_i;
  wire irq_pending_i;
  input irq_pending_i_t0;
  wire irq_pending_i_t0;
  input [17:0] irqs_i;
  wire [17:0] irqs_i;
  input [17:0] irqs_i_t0;
  wire [17:0] irqs_i_t0;
  wire jump_in_dec;
  wire jump_in_dec_t0;
  wire jump_set;
  wire jump_set_dec;
  wire jump_set_dec_t0;
  wire jump_set_raw;
  wire jump_set_raw_t0;
  wire jump_set_t0;
  input lsu_addr_incr_req_i;
  wire lsu_addr_incr_req_i;
  input lsu_addr_incr_req_i_t0;
  wire lsu_addr_incr_req_i_t0;
  input [31:0] lsu_addr_last_i;
  wire [31:0] lsu_addr_last_i;
  input [31:0] lsu_addr_last_i_t0;
  wire [31:0] lsu_addr_last_i_t0;
  input lsu_load_err_i;
  wire lsu_load_err_i;
  input lsu_load_err_i_t0;
  wire lsu_load_err_i_t0;
  wire lsu_req_dec;
  wire lsu_req_dec_t0;
  input lsu_req_done_i;
  wire lsu_req_done_i;
  input lsu_req_done_i_t0;
  wire lsu_req_done_i_t0;
  output lsu_req_o;
  wire lsu_req_o;
  output lsu_req_o_t0;
  wire lsu_req_o_t0;
  input lsu_resp_valid_i;
  wire lsu_resp_valid_i;
  input lsu_resp_valid_i_t0;
  wire lsu_resp_valid_i_t0;
  output lsu_sign_ext_o;
  wire lsu_sign_ext_o;
  output lsu_sign_ext_o_t0;
  wire lsu_sign_ext_o_t0;
  input lsu_store_err_i;
  wire lsu_store_err_i;
  input lsu_store_err_i_t0;
  wire lsu_store_err_i_t0;
  output [1:0] lsu_type_o;
  wire [1:0] lsu_type_o;
  output [1:0] lsu_type_o_t0;
  wire [1:0] lsu_type_o_t0;
  output [31:0] lsu_wdata_o;
  wire [31:0] lsu_wdata_o;
  output [31:0] lsu_wdata_o_t0;
  wire [31:0] lsu_wdata_o_t0;
  output lsu_we_o;
  wire lsu_we_o;
  output lsu_we_o_t0;
  wire lsu_we_o_t0;
  wire mret_insn_dec;
  wire mret_insn_dec_t0;
  wire mult_en_dec;
  wire mult_en_dec_t0;
  output mult_en_ex_o;
  wire mult_en_ex_o;
  output mult_en_ex_o_t0;
  wire mult_en_ex_o_t0;
  output mult_sel_ex_o;
  wire mult_sel_ex_o;
  output mult_sel_ex_o_t0;
  wire mult_sel_ex_o_t0;
  wire multdiv_en_dec;
  wire multdiv_en_dec_t0;
  output [31:0] multdiv_operand_a_ex_o;
  wire [31:0] multdiv_operand_a_ex_o;
  output [31:0] multdiv_operand_a_ex_o_t0;
  wire [31:0] multdiv_operand_a_ex_o_t0;
  output [31:0] multdiv_operand_b_ex_o;
  wire [31:0] multdiv_operand_b_ex_o;
  output [31:0] multdiv_operand_b_ex_o_t0;
  wire [31:0] multdiv_operand_b_ex_o_t0;
  output [1:0] multdiv_operator_ex_o;
  wire [1:0] multdiv_operator_ex_o;
  output [1:0] multdiv_operator_ex_o_t0;
  wire [1:0] multdiv_operator_ex_o_t0;
  output multdiv_ready_id_o;
  wire multdiv_ready_id_o;
  output multdiv_ready_id_o_t0;
  wire multdiv_ready_id_o_t0;
  output [1:0] multdiv_signed_mode_ex_o;
  wire [1:0] multdiv_signed_mode_ex_o;
  output [1:0] multdiv_signed_mode_ex_o_t0;
  wire [1:0] multdiv_signed_mode_ex_o_t0;
  wire multicycle_done;
  wire multicycle_done_t0;
  output nmi_mode_o;
  wire nmi_mode_o;
  output nmi_mode_o_t0;
  wire nmi_mode_o_t0;
  output nt_branch_mispredict_o;
  wire nt_branch_mispredict_o;
  output nt_branch_mispredict_o_t0;
  wire nt_branch_mispredict_o_t0;
  input outstanding_load_wb_i;
  wire outstanding_load_wb_i;
  input outstanding_load_wb_i_t0;
  wire outstanding_load_wb_i_t0;
  input outstanding_store_wb_i;
  wire outstanding_store_wb_i;
  input outstanding_store_wb_i_t0;
  wire outstanding_store_wb_i_t0;
  input [31:0] pc_id_i;
  wire [31:0] pc_id_i;
  input [31:0] pc_id_i_t0;
  wire [31:0] pc_id_i_t0;
  output [2:0] pc_mux_o;
  wire [2:0] pc_mux_o;
  output [2:0] pc_mux_o_t0;
  wire [2:0] pc_mux_o_t0;
  output pc_set_o;
  wire pc_set_o;
  output pc_set_o_t0;
  wire pc_set_o_t0;
  output pc_set_spec_o;
  wire pc_set_spec_o;
  output pc_set_spec_o_t0;
  wire pc_set_spec_o_t0;
  output perf_branch_o;
  wire perf_branch_o;
  output perf_branch_o_t0;
  wire perf_branch_o_t0;
  output perf_div_wait_o;
  wire perf_div_wait_o;
  output perf_div_wait_o_t0;
  wire perf_div_wait_o_t0;
  output perf_dside_wait_o;
  wire perf_dside_wait_o;
  output perf_dside_wait_o_t0;
  wire perf_dside_wait_o_t0;
  output perf_jump_o;
  wire perf_jump_o;
  output perf_jump_o_t0;
  wire perf_jump_o_t0;
  output perf_mul_wait_o;
  wire perf_mul_wait_o;
  output perf_mul_wait_o_t0;
  wire perf_mul_wait_o_t0;
  output perf_tbranch_o;
  wire perf_tbranch_o;
  output perf_tbranch_o_t0;
  wire perf_tbranch_o_t0;
  input [1:0] priv_mode_i;
  wire [1:0] priv_mode_i;
  input [1:0] priv_mode_i_t0;
  wire [1:0] priv_mode_i_t0;
  input ready_wb_i;
  wire ready_wb_i;
  input ready_wb_i_t0;
  wire ready_wb_i_t0;
  input [31:0] result_ex_i;
  wire [31:0] result_ex_i;
  input [31:0] result_ex_i_t0;
  wire [31:0] result_ex_i_t0;
  output [4:0] rf_raddr_a_o;
  wire [4:0] rf_raddr_a_o;
  output [4:0] rf_raddr_a_o_t0;
  wire [4:0] rf_raddr_a_o_t0;
  output [4:0] rf_raddr_b_o;
  wire [4:0] rf_raddr_b_o;
  output [4:0] rf_raddr_b_o_t0;
  wire [4:0] rf_raddr_b_o_t0;
  output rf_rd_a_wb_match_o;
  wire rf_rd_a_wb_match_o;
  output rf_rd_a_wb_match_o_t0;
  wire rf_rd_a_wb_match_o_t0;
  output rf_rd_b_wb_match_o;
  wire rf_rd_b_wb_match_o;
  output rf_rd_b_wb_match_o_t0;
  wire rf_rd_b_wb_match_o_t0;
  input [31:0] rf_rdata_a_i;
  wire [31:0] rf_rdata_a_i;
  input [31:0] rf_rdata_a_i_t0;
  wire [31:0] rf_rdata_a_i_t0;
  input [31:0] rf_rdata_b_i;
  wire [31:0] rf_rdata_b_i;
  input [31:0] rf_rdata_b_i_t0;
  wire [31:0] rf_rdata_b_i_t0;
  wire rf_ren_a_dec;
  wire rf_ren_a_dec_t0;
  output rf_ren_a_o;
  wire rf_ren_a_o;
  output rf_ren_a_o_t0;
  wire rf_ren_a_o_t0;
  wire rf_ren_b_dec;
  wire rf_ren_b_dec_t0;
  output rf_ren_b_o;
  wire rf_ren_b_o;
  output rf_ren_b_o_t0;
  wire rf_ren_b_o_t0;
  output [4:0] rf_waddr_id_o;
  wire [4:0] rf_waddr_id_o;
  output [4:0] rf_waddr_id_o_t0;
  wire [4:0] rf_waddr_id_o_t0;
  input [4:0] rf_waddr_wb_i;
  wire [4:0] rf_waddr_wb_i;
  input [4:0] rf_waddr_wb_i_t0;
  wire [4:0] rf_waddr_wb_i_t0;
  input [31:0] rf_wdata_fwd_wb_i;
  wire [31:0] rf_wdata_fwd_wb_i;
  input [31:0] rf_wdata_fwd_wb_i_t0;
  wire [31:0] rf_wdata_fwd_wb_i_t0;
  output [31:0] rf_wdata_id_o;
  wire [31:0] rf_wdata_id_o;
  output [31:0] rf_wdata_id_o_t0;
  wire [31:0] rf_wdata_id_o_t0;
  wire rf_wdata_sel;
  wire rf_wdata_sel_t0;
  wire rf_we_dec;
  wire rf_we_dec_t0;
  output rf_we_id_o;
  wire rf_we_id_o;
  output rf_we_id_o_t0;
  wire rf_we_id_o_t0;
  wire rf_we_raw;
  wire rf_we_raw_t0;
  input rf_write_wb_i;
  wire rf_write_wb_i;
  input rf_write_wb_i_t0;
  wire rf_write_wb_i_t0;
  input rst_ni;
  wire rst_ni;
  wire stall_alu;
  wire stall_alu_t0;
  wire stall_branch;
  wire stall_branch_t0;
  wire stall_id;
  wire stall_id_t0;
  wire stall_jump;
  wire stall_jump_t0;
  wire stall_ld_hz;
  wire stall_ld_hz_t0;
  wire stall_mem;
  wire stall_mem_t0;
  wire stall_multdiv;
  wire stall_multdiv_t0;
  wire stall_wb;
  wire stall_wb_t0;
  input trigger_match_i;
  wire trigger_match_i;
  input trigger_match_i_t0;
  wire trigger_match_i_t0;
  wire wb_exception;
  wire wb_exception_t0;
  wire wfi_insn_dec;
  wire wfi_insn_dec_t0;
  wire [31:0] zimm_rs1_type;
  wire [31:0] zimm_rs1_type_t0;
  assign rf_ren_a_o = _0060_ & rf_ren_a_dec;
  assign _0060_ = _0058_ & _0944_;
  assign rf_ren_b_o = _0060_ & rf_ren_b_dec;
  assign _0062_ = rf_we_raw & instr_executing;
  assign rf_we_id_o = _0062_ & _0129_;
  assign illegal_insn_o = instr_valid_i & _0954_;
  assign _0064_ = data_req_allowed & lsu_req_dec;
  assign _0066_ = csr_access_o & instr_executing;
  assign csr_op_en_o = _0066_ & instr_id_done_o;
  assign branch_jump_set_done_d = _0958_ & _0945_;
  assign jump_set = jump_set_raw & _0135_;
  assign branch_set = branch_set_raw & _0135_;
  assign branch_set_spec = branch_set_raw_spec & _0135_;
  assign _0068_ = rf_we_dec & ex_valid_i;
  assign _0070_ = multicycle_done & ready_wb_i;
  assign _0071_ = _0946_ & _0947_;
  assign en_wb_o = _0071_ & instr_executing;
  assign instr_first_cycle_id_o = instr_valid_i & _0109_;
  assign \gen_stall_mem.outstanding_memory_access  = _0969_ & _0948_;
  assign _0058_ = instr_valid_i & _0150_;
  assign _0073_ = _0058_ & controller_run;
  assign instr_executing_spec = _0073_ & _0138_;
  assign _0077_ = _0075_ & _0138_;
  assign instr_executing = _0077_ & data_req_allowed;
  assign _0079_ = lsu_req_dec & _0162_;
  assign stall_mem = instr_valid_i & _0973_;
  assign rf_rd_a_wb_match_o = _0926_ & _1027_;
  assign rf_rd_b_wb_match_o = _0928_ & _1029_;
  assign \gen_stall_mem.rf_rd_a_hz  = rf_rd_a_wb_match_o & rf_ren_a_o;
  assign \gen_stall_mem.rf_rd_b_hz  = rf_rd_b_wb_match_o & rf_ren_b_o;
  assign _0081_ = rf_rd_a_wb_match_o & rf_write_wb_i;
  assign _0083_ = rf_rd_b_wb_match_o & rf_write_wb_i;
  assign stall_ld_hz = outstanding_load_wb_i & _0975_;
  assign instr_id_done_o = en_wb_o & ready_wb_i;
  assign stall_wb = en_wb_o & _0951_;
  assign _0075_ = instr_valid_i & _0950_;
  assign perf_dside_wait_o = _0075_ & _0977_;
  assign _0085_ = _0952_ & _0953_;
  assign _0087_ = _0085_ & _0128_;
  assign _0089_ = _0087_ & _0129_;
  assign instr_perf_count_id_o = _0089_ & _0150_;
  assign perf_mul_wait_o = stall_multdiv & mult_en_dec;
  assign perf_div_wait_o = stall_multdiv & div_en_dec;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) branch_jump_set_done_q_t0 <= 1'h0;
    else branch_jump_set_done_q_t0 <= branch_jump_set_done_d_t0;
  assign _0093_ = ~ _0091_;
  assign _0094_ = ~ imd_val_we_ex_i[1];
  assign _0095_ = ~ imd_val_we_ex_i[0];
  assign _0825_ = _0006_ ^ id_fsm_q;
  assign _0826_ = imd_val_d_ex_i[33:0] ^ imd_val_q_ex_o[33:0];
  assign _0827_ = imd_val_d_ex_i[67:34] ^ imd_val_q_ex_o[67:34];
  assign _0686_ = _0007_ | id_fsm_q_t0;
  assign _0690_ = imd_val_d_ex_i_t0[33:0] | imd_val_q_ex_o_t0[33:0];
  assign _0694_ = imd_val_d_ex_i_t0[67:34] | imd_val_q_ex_o_t0[67:34];
  assign _0687_ = _0825_ | _0686_;
  assign _0691_ = _0826_ | _0690_;
  assign _0695_ = _0827_ | _0694_;
  assign _0328_ = _0091_ & _0007_;
  assign _0331_ = { imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1] } & imd_val_d_ex_i_t0[33:0];
  assign _0334_ = { imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0] } & imd_val_d_ex_i_t0[67:34];
  assign _0329_ = _0093_ & id_fsm_q_t0;
  assign _0332_ = { _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_ } & imd_val_q_ex_o_t0[33:0];
  assign _0335_ = { _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_ } & imd_val_q_ex_o_t0[67:34];
  assign _0330_ = _0687_ & _0092_;
  assign _0333_ = _0691_ & { imd_val_we_ex_i_t0[1], imd_val_we_ex_i_t0[1], imd_val_we_ex_i_t0[1], imd_val_we_ex_i_t0[1], imd_val_we_ex_i_t0[1], imd_val_we_ex_i_t0[1], imd_val_we_ex_i_t0[1], imd_val_we_ex_i_t0[1], imd_val_we_ex_i_t0[1], imd_val_we_ex_i_t0[1], imd_val_we_ex_i_t0[1], imd_val_we_ex_i_t0[1], imd_val_we_ex_i_t0[1], imd_val_we_ex_i_t0[1], imd_val_we_ex_i_t0[1], imd_val_we_ex_i_t0[1], imd_val_we_ex_i_t0[1], imd_val_we_ex_i_t0[1], imd_val_we_ex_i_t0[1], imd_val_we_ex_i_t0[1], imd_val_we_ex_i_t0[1], imd_val_we_ex_i_t0[1], imd_val_we_ex_i_t0[1], imd_val_we_ex_i_t0[1], imd_val_we_ex_i_t0[1], imd_val_we_ex_i_t0[1], imd_val_we_ex_i_t0[1], imd_val_we_ex_i_t0[1], imd_val_we_ex_i_t0[1], imd_val_we_ex_i_t0[1], imd_val_we_ex_i_t0[1], imd_val_we_ex_i_t0[1], imd_val_we_ex_i_t0[1], imd_val_we_ex_i_t0[1] };
  assign _0336_ = _0695_ & { imd_val_we_ex_i_t0[0], imd_val_we_ex_i_t0[0], imd_val_we_ex_i_t0[0], imd_val_we_ex_i_t0[0], imd_val_we_ex_i_t0[0], imd_val_we_ex_i_t0[0], imd_val_we_ex_i_t0[0], imd_val_we_ex_i_t0[0], imd_val_we_ex_i_t0[0], imd_val_we_ex_i_t0[0], imd_val_we_ex_i_t0[0], imd_val_we_ex_i_t0[0], imd_val_we_ex_i_t0[0], imd_val_we_ex_i_t0[0], imd_val_we_ex_i_t0[0], imd_val_we_ex_i_t0[0], imd_val_we_ex_i_t0[0], imd_val_we_ex_i_t0[0], imd_val_we_ex_i_t0[0], imd_val_we_ex_i_t0[0], imd_val_we_ex_i_t0[0], imd_val_we_ex_i_t0[0], imd_val_we_ex_i_t0[0], imd_val_we_ex_i_t0[0], imd_val_we_ex_i_t0[0], imd_val_we_ex_i_t0[0], imd_val_we_ex_i_t0[0], imd_val_we_ex_i_t0[0], imd_val_we_ex_i_t0[0], imd_val_we_ex_i_t0[0], imd_val_we_ex_i_t0[0], imd_val_we_ex_i_t0[0], imd_val_we_ex_i_t0[0], imd_val_we_ex_i_t0[0] };
  assign _0688_ = _0328_ | _0329_;
  assign _0692_ = _0331_ | _0332_;
  assign _0696_ = _0334_ | _0335_;
  assign _0689_ = _0688_ | _0330_;
  assign _0693_ = _0692_ | _0333_;
  assign _0697_ = _0696_ | _0336_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) id_fsm_q_t0 <= 1'h0;
    else id_fsm_q_t0 <= _0689_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) imd_val_q_ex_o_t0[33:0] <= 34'h000000000;
    else imd_val_q_ex_o_t0[33:0] <= _0693_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) imd_val_q_ex_o_t0[67:34] <= 34'h000000000;
    else imd_val_q_ex_o_t0[67:34] <= _0697_;
  assign _0201_ = _0061_ & rf_ren_a_dec;
  assign _0204_ = _0059_ & _0944_;
  assign _0207_ = _0061_ & rf_ren_b_dec;
  assign _0210_ = rf_we_raw_t0 & instr_executing;
  assign _0213_ = _0063_ & _0129_;
  assign _0216_ = instr_valid_i_t0 & _0954_;
  assign _0219_ = data_req_allowed_t0 & lsu_req_dec;
  assign _0222_ = csr_access_o_t0 & instr_executing;
  assign _0225_ = _0067_ & instr_id_done_o;
  assign _0228_ = _0959_ & _0945_;
  assign _0231_ = jump_set_raw_t0 & _0135_;
  assign _0234_ = branch_set_raw_t0 & _0135_;
  assign _0237_ = branch_set_raw_spec_t0 & _0135_;
  assign _0240_ = rf_we_dec_t0 & ex_valid_i;
  assign _0243_ = multicycle_done_t0 & ready_wb_i;
  assign _0246_ = stall_id_t0 & _0947_;
  assign _0249_ = _0072_ & instr_executing;
  assign _0252_ = instr_valid_i_t0 & _0109_;
  assign _0255_ = _0970_ & _0948_;
  assign _0258_ = instr_valid_i_t0 & _0150_;
  assign _0261_ = _0059_ & controller_run;
  assign _0264_ = _0074_ & _0138_;
  assign _0267_ = _0076_ & _0138_;
  assign _0270_ = _0078_ & data_req_allowed;
  assign _0273_ = lsu_req_dec_t0 & _0162_;
  assign _0276_ = instr_valid_i_t0 & _0973_;
  assign _0279_ = _0927_ & _1027_;
  assign _0282_ = _0929_ & _1029_;
  assign _0285_ = rf_rd_a_wb_match_o_t0 & rf_ren_a_o;
  assign _0288_ = rf_rd_b_wb_match_o_t0 & rf_ren_b_o;
  assign _0291_ = rf_rd_a_wb_match_o_t0 & rf_write_wb_i;
  assign _0294_ = rf_rd_b_wb_match_o_t0 & rf_write_wb_i;
  assign _0297_ = outstanding_load_wb_i_t0 & _0975_;
  assign _0300_ = en_wb_o_t0 & ready_wb_i;
  assign _0303_ = en_wb_o_t0 & _0951_;
  assign _0304_ = instr_valid_i_t0 & _0950_;
  assign _0307_ = _0076_ & _0977_;
  assign _0310_ = ebrk_insn_t0 & _0953_;
  assign _0313_ = _0086_ & _0128_;
  assign _0316_ = _0088_ & _0129_;
  assign _0319_ = _0090_ & _0150_;
  assign _0322_ = stall_multdiv_t0 & mult_en_dec;
  assign _0325_ = stall_multdiv_t0 & div_en_dec;
  assign _0202_ = rf_ren_a_dec_t0 & _0060_;
  assign _0205_ = illegal_insn_o_t0 & _0058_;
  assign _0208_ = rf_ren_b_dec_t0 & _0060_;
  assign _0211_ = instr_executing_t0 & rf_we_raw;
  assign _0214_ = illegal_csr_insn_i_t0 & _0062_;
  assign _0217_ = _0955_ & instr_valid_i;
  assign _0220_ = lsu_req_dec_t0 & data_req_allowed;
  assign _0223_ = instr_executing_t0 & csr_access_o;
  assign _0226_ = instr_id_done_o_t0 & _0066_;
  assign _0229_ = instr_valid_clear_o_t0 & _0958_;
  assign _0232_ = branch_jump_set_done_q_t0 & jump_set_raw;
  assign _0235_ = branch_jump_set_done_q_t0 & branch_set_raw;
  assign _0238_ = branch_jump_set_done_q_t0 & branch_set_raw_spec;
  assign _0244_ = ready_wb_i_t0 & multicycle_done;
  assign _0247_ = flush_id_t0 & _0946_;
  assign _0250_ = instr_executing_t0 & _0071_;
  assign _0253_ = id_fsm_q_t0 & instr_valid_i;
  assign _0256_ = lsu_resp_valid_i_t0 & _0969_;
  assign _0259_ = instr_fetch_err_i_t0 & instr_valid_i;
  assign _0262_ = controller_run_t0 & _0058_;
  assign _0265_ = stall_ld_hz_t0 & _0073_;
  assign _0268_ = stall_ld_hz_t0 & _0075_;
  assign _0271_ = data_req_allowed_t0 & _0077_;
  assign _0274_ = lsu_req_done_i_t0 & lsu_req_dec;
  assign _0277_ = _0974_ & instr_valid_i;
  assign _0280_ = _1028_ & _0926_;
  assign _0283_ = _1030_ & _0928_;
  assign _0286_ = rf_ren_a_o_t0 & rf_rd_a_wb_match_o;
  assign _0289_ = rf_ren_b_o_t0 & rf_rd_b_wb_match_o;
  assign _0292_ = rf_write_wb_i_t0 & rf_rd_a_wb_match_o;
  assign _0295_ = rf_write_wb_i_t0 & rf_rd_b_wb_match_o;
  assign _0298_ = _0976_ & outstanding_load_wb_i;
  assign _0301_ = ready_wb_i_t0 & en_wb_o;
  assign _0305_ = \gen_stall_mem.instr_kill_t0  & instr_valid_i;
  assign _0308_ = _0978_ & _0075_;
  assign _0311_ = ecall_insn_dec_t0 & _0952_;
  assign _0314_ = illegal_insn_dec_t0 & _0085_;
  assign _0317_ = illegal_csr_insn_i_t0 & _0087_;
  assign _0320_ = instr_fetch_err_i_t0 & _0089_;
  assign _0323_ = mult_en_dec_t0 & stall_multdiv;
  assign _0326_ = div_en_dec_t0 & stall_multdiv;
  assign _0203_ = _0061_ & rf_ren_a_dec_t0;
  assign _0206_ = _0059_ & illegal_insn_o_t0;
  assign _0209_ = _0061_ & rf_ren_b_dec_t0;
  assign _0212_ = rf_we_raw_t0 & instr_executing_t0;
  assign _0215_ = _0063_ & illegal_csr_insn_i_t0;
  assign _0218_ = instr_valid_i_t0 & _0955_;
  assign _0221_ = data_req_allowed_t0 & lsu_req_dec_t0;
  assign _0224_ = csr_access_o_t0 & instr_executing_t0;
  assign _0227_ = _0067_ & instr_id_done_o_t0;
  assign _0230_ = _0959_ & instr_valid_clear_o_t0;
  assign _0233_ = jump_set_raw_t0 & branch_jump_set_done_q_t0;
  assign _0236_ = branch_set_raw_t0 & branch_jump_set_done_q_t0;
  assign _0239_ = branch_set_raw_spec_t0 & branch_jump_set_done_q_t0;
  assign _0242_ = rf_we_dec_t0 & ex_valid_i_t0;
  assign _0245_ = multicycle_done_t0 & ready_wb_i_t0;
  assign _0248_ = stall_id_t0 & flush_id_t0;
  assign _0251_ = _0072_ & instr_executing_t0;
  assign _0254_ = instr_valid_i_t0 & id_fsm_q_t0;
  assign _0257_ = _0970_ & lsu_resp_valid_i_t0;
  assign _0260_ = instr_valid_i_t0 & instr_fetch_err_i_t0;
  assign _0263_ = _0059_ & controller_run_t0;
  assign _0266_ = _0074_ & stall_ld_hz_t0;
  assign _0269_ = _0076_ & stall_ld_hz_t0;
  assign _0272_ = _0078_ & data_req_allowed_t0;
  assign _0275_ = lsu_req_dec_t0 & lsu_req_done_i_t0;
  assign _0278_ = instr_valid_i_t0 & _0974_;
  assign _0281_ = _0927_ & _1028_;
  assign _0284_ = _0929_ & _1030_;
  assign _0287_ = rf_rd_a_wb_match_o_t0 & rf_ren_a_o_t0;
  assign _0290_ = rf_rd_b_wb_match_o_t0 & rf_ren_b_o_t0;
  assign _0293_ = rf_rd_a_wb_match_o_t0 & rf_write_wb_i_t0;
  assign _0296_ = rf_rd_b_wb_match_o_t0 & rf_write_wb_i_t0;
  assign _0299_ = outstanding_load_wb_i_t0 & _0976_;
  assign _0302_ = en_wb_o_t0 & ready_wb_i_t0;
  assign _0306_ = instr_valid_i_t0 & \gen_stall_mem.instr_kill_t0 ;
  assign _0309_ = _0076_ & _0978_;
  assign _0312_ = ebrk_insn_t0 & ecall_insn_dec_t0;
  assign _0315_ = _0086_ & illegal_insn_dec_t0;
  assign _0318_ = _0088_ & illegal_csr_insn_i_t0;
  assign _0321_ = _0090_ & instr_fetch_err_i_t0;
  assign _0324_ = stall_multdiv_t0 & mult_en_dec_t0;
  assign _0327_ = stall_multdiv_t0 & div_en_dec_t0;
  assign _0643_ = _0201_ | _0202_;
  assign _0644_ = _0204_ | _0205_;
  assign _0645_ = _0207_ | _0208_;
  assign _0646_ = _0210_ | _0211_;
  assign _0647_ = _0213_ | _0214_;
  assign _0648_ = _0216_ | _0217_;
  assign _0649_ = _0219_ | _0220_;
  assign _0650_ = _0222_ | _0223_;
  assign _0651_ = _0225_ | _0226_;
  assign _0652_ = _0228_ | _0229_;
  assign _0653_ = _0231_ | _0232_;
  assign _0654_ = _0234_ | _0235_;
  assign _0655_ = _0237_ | _0238_;
  assign _0656_ = _0240_ | _0241_;
  assign _0657_ = _0243_ | _0244_;
  assign _0658_ = _0246_ | _0247_;
  assign _0659_ = _0249_ | _0250_;
  assign _0660_ = _0252_ | _0253_;
  assign _0661_ = _0255_ | _0256_;
  assign _0662_ = _0258_ | _0259_;
  assign _0663_ = _0261_ | _0262_;
  assign _0664_ = _0264_ | _0265_;
  assign _0665_ = _0267_ | _0268_;
  assign _0666_ = _0270_ | _0271_;
  assign _0667_ = _0273_ | _0274_;
  assign _0668_ = _0276_ | _0277_;
  assign _0669_ = _0279_ | _0280_;
  assign _0670_ = _0282_ | _0283_;
  assign _0671_ = _0285_ | _0286_;
  assign _0672_ = _0288_ | _0289_;
  assign _0673_ = _0291_ | _0292_;
  assign _0674_ = _0294_ | _0295_;
  assign _0675_ = _0297_ | _0298_;
  assign _0676_ = _0300_ | _0301_;
  assign _0677_ = _0303_ | _0301_;
  assign _0678_ = _0304_ | _0305_;
  assign _0679_ = _0307_ | _0308_;
  assign _0680_ = _0310_ | _0311_;
  assign _0681_ = _0313_ | _0314_;
  assign _0682_ = _0316_ | _0317_;
  assign _0683_ = _0319_ | _0320_;
  assign _0684_ = _0322_ | _0323_;
  assign _0685_ = _0325_ | _0326_;
  assign rf_ren_a_o_t0 = _0643_ | _0203_;
  assign _0061_ = _0644_ | _0206_;
  assign rf_ren_b_o_t0 = _0645_ | _0209_;
  assign _0063_ = _0646_ | _0212_;
  assign rf_we_id_o_t0 = _0647_ | _0215_;
  assign illegal_insn_o_t0 = _0648_ | _0218_;
  assign _0065_ = _0649_ | _0221_;
  assign _0067_ = _0650_ | _0224_;
  assign csr_op_en_o_t0 = _0651_ | _0227_;
  assign branch_jump_set_done_d_t0 = _0652_ | _0230_;
  assign jump_set_t0 = _0653_ | _0233_;
  assign branch_set_t0 = _0654_ | _0236_;
  assign branch_set_spec_t0 = _0655_ | _0239_;
  assign _0069_ = _0656_ | _0242_;
  assign _0057_ = _0657_ | _0245_;
  assign _0072_ = _0658_ | _0248_;
  assign en_wb_o_t0 = _0659_ | _0251_;
  assign instr_first_cycle_id_o_t0 = _0660_ | _0254_;
  assign data_req_allowed_t0 = _0661_ | _0257_;
  assign _0059_ = _0662_ | _0260_;
  assign _0074_ = _0663_ | _0263_;
  assign instr_executing_spec_t0 = _0664_ | _0266_;
  assign _0078_ = _0665_ | _0269_;
  assign instr_executing_t0 = _0666_ | _0272_;
  assign _0080_ = _0667_ | _0275_;
  assign stall_mem_t0 = _0668_ | _0278_;
  assign rf_rd_a_wb_match_o_t0 = _0669_ | _0281_;
  assign rf_rd_b_wb_match_o_t0 = _0670_ | _0284_;
  assign \gen_stall_mem.rf_rd_a_hz_t0  = _0671_ | _0287_;
  assign \gen_stall_mem.rf_rd_b_hz_t0  = _0672_ | _0290_;
  assign _0082_ = _0673_ | _0293_;
  assign _0084_ = _0674_ | _0296_;
  assign stall_ld_hz_t0 = _0675_ | _0299_;
  assign instr_id_done_o_t0 = _0676_ | _0302_;
  assign stall_wb_t0 = _0677_ | _0302_;
  assign _0076_ = _0678_ | _0306_;
  assign perf_dside_wait_o_t0 = _0679_ | _0309_;
  assign _0086_ = _0680_ | _0312_;
  assign _0088_ = _0681_ | _0315_;
  assign _0090_ = _0682_ | _0318_;
  assign instr_perf_count_id_o_t0 = _0683_ | _0321_;
  assign perf_mul_wait_o_t0 = _0684_ | _0324_;
  assign perf_div_wait_o_t0 = _0685_ | _0327_;
  assign _0186_ = | instr_rdata_i_t0[31:20];
  assign _0187_ = | { rf_waddr_wb_i_t0, rf_raddr_a_o_t0 };
  assign _0188_ = | { rf_waddr_wb_i_t0, rf_raddr_b_o_t0 };
  assign _0192_ = | alu_op_a_mux_sel_t0;
  assign _0741_ = rf_waddr_wb_i_t0 | rf_raddr_a_o_t0;
  assign _0742_ = rf_waddr_wb_i_t0 | rf_raddr_b_o_t0;
  assign _0114_ = ~ csr_op_o_t0;
  assign _0115_ = ~ instr_rdata_i_t0[31:20];
  assign _0116_ = ~ _0741_;
  assign _0117_ = ~ _0742_;
  assign _0156_ = ~ imm_b_mux_sel_t0;
  assign _0157_ = ~ bt_b_mux_sel_t0;
  assign _0169_ = ~ alu_op_a_mux_sel_t0;
  assign _0403_ = csr_op_o & _0114_;
  assign _0406_ = instr_rdata_i[31:20] & _0115_;
  assign _0413_ = rf_waddr_wb_i & _0116_;
  assign _0415_ = rf_waddr_wb_i & _0117_;
  assign _0486_ = imm_b_mux_sel & _0156_;
  assign _0490_ = bt_b_mux_sel & _0157_;
  assign _0593_ = alu_op_a_mux_sel & _0169_;
  assign _0404_ = 2'h1 & _0114_;
  assign _0405_ = 2'h2 & _0114_;
  assign _0407_ = 12'h300 & _0115_;
  assign _0408_ = 12'h304 & _0115_;
  assign _0409_ = 12'h7b0 & _0115_;
  assign _0410_ = 12'h7b1 & _0115_;
  assign _0411_ = 12'h7b2 & _0115_;
  assign _0412_ = 12'h7b3 & _0115_;
  assign _0414_ = rf_raddr_a_o & _0116_;
  assign _0416_ = rf_raddr_b_o & _0117_;
  assign _0487_ = 3'h5 & _0156_;
  assign _0488_ = 3'h3 & _0156_;
  assign _0489_ = 3'h1 & _0156_;
  assign _0491_ = 3'h4 & _0157_;
  assign _0492_ = 3'h2 & _0157_;
  assign _0594_ = 2'h3 & _0169_;
  assign _0595_ = 2'h2 & _0169_;
  assign _0596_ = 2'h1 & _0169_;
  assign _0878_ = _0403_ == _0404_;
  assign _0879_ = _0403_ == _0405_;
  assign _0880_ = _0406_ == _0407_;
  assign _0881_ = _0406_ == _0408_;
  assign _0882_ = _0406_ == _0409_;
  assign _0883_ = _0406_ == _0410_;
  assign _0884_ = _0406_ == _0411_;
  assign _0885_ = _0406_ == _0412_;
  assign _0886_ = _0413_ == _0414_;
  assign _0887_ = _0415_ == _0416_;
  assign _0888_ = _0486_ == _0487_;
  assign _0889_ = _0486_ == _0488_;
  assign _0890_ = _0486_ == _0489_;
  assign _0891_ = _0490_ == _0491_;
  assign _0892_ = _0490_ == _0492_;
  assign _0893_ = _0593_ == _0594_;
  assign _0894_ = _0593_ == _0595_;
  assign _0895_ = _0593_ == _0596_;
  assign _0911_ = _0878_ & _0185_;
  assign _0913_ = _0879_ & _0185_;
  assign _0915_ = _0880_ & _0186_;
  assign _0917_ = _0881_ & _0186_;
  assign _0919_ = _0882_ & _0186_;
  assign _0921_ = _0883_ & _0186_;
  assign _0923_ = _0884_ & _0186_;
  assign _0925_ = _0885_ & _0186_;
  assign _0927_ = _0886_ & _0187_;
  assign _0929_ = _0887_ & _0188_;
  assign _0980_ = _0888_ & _0189_;
  assign _0982_ = _0889_ & _0189_;
  assign _0984_ = _0890_ & _0189_;
  assign _0988_ = _0891_ & _0190_;
  assign _0990_ = _0892_ & _0190_;
  assign _1022_ = _0893_ & _0192_;
  assign _1024_ = _0894_ & _0192_;
  assign _1026_ = _0895_ & _0192_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) id_fsm_q <= 1'h0;
    else if (_0091_) id_fsm_q <= _0006_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) imd_val_q_ex_o[33:0] <= 34'h000000000;
    else if (imd_val_we_ex_i[1]) imd_val_q_ex_o[33:0] <= imd_val_d_ex_i[33:0];
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) imd_val_q_ex_o[67:34] <= 34'h000000000;
    else if (imd_val_we_ex_i[0]) imd_val_q_ex_o[67:34] <= imd_val_d_ex_i[67:34];
  assign _0417_ = csr_op_en_o_t0 & _0934_;
  assign _0420_ = csr_op_en_o_t0 & _0942_;
  assign _0418_ = _0935_ & csr_op_en_o;
  assign _0421_ = _0943_ & csr_op_en_o;
  assign _0419_ = csr_op_en_o_t0 & _0935_;
  assign _0422_ = csr_op_en_o_t0 & _0943_;
  assign _0743_ = _0417_ | _0418_;
  assign _0744_ = _0420_ | _0421_;
  assign _0931_ = _0743_ | _0419_;
  assign _0933_ = _0744_ | _0422_;
  assign _0185_ = | csr_op_o_t0;
  assign _0189_ = | imm_b_mux_sel_t0;
  assign _0190_ = | bt_b_mux_sel_t0;
  assign _0191_ = | bt_a_mux_sel_t0;
  assign _0193_ = | rf_raddr_a_o_t0;
  assign _0194_ = | rf_raddr_b_o_t0;
  assign _0159_ = ~ bt_a_mux_sel_t0;
  assign _0170_ = ~ rf_raddr_a_o_t0;
  assign _0171_ = ~ rf_raddr_b_o_t0;
  assign _0496_ = bt_a_mux_sel & _0159_;
  assign _0597_ = rf_raddr_a_o & _0170_;
  assign _0598_ = rf_raddr_b_o & _0171_;
  assign _0195_ = ! _0403_;
  assign _0196_ = ! _0486_;
  assign _0197_ = ! _0490_;
  assign _0198_ = ! _0496_;
  assign _0199_ = ! _0597_;
  assign _0200_ = ! _0598_;
  assign _0943_ = _0195_ & _0185_;
  assign _0986_ = _0196_ & _0189_;
  assign _0992_ = _0197_ & _0190_;
  assign _0994_ = _0198_ & _0191_;
  assign _1028_ = _0199_ & _0193_;
  assign _1030_ = _0200_ & _0194_;
  assign _0118_ = ~ _0910_;
  assign _0120_ = ~ _0914_;
  assign _0122_ = ~ _0918_;
  assign _0124_ = ~ _0937_;
  assign _0126_ = ~ _0939_;
  assign _0119_ = ~ _0912_;
  assign _0121_ = ~ _0916_;
  assign _0123_ = ~ _0920_;
  assign _0125_ = ~ _0922_;
  assign _0127_ = ~ _0924_;
  assign _0423_ = _0911_ & _0119_;
  assign _0426_ = _0915_ & _0121_;
  assign _0429_ = _0919_ & _0123_;
  assign _0432_ = _0938_ & _0125_;
  assign _0435_ = _0940_ & _0127_;
  assign _0424_ = _0913_ & _0118_;
  assign _0427_ = _0917_ & _0120_;
  assign _0430_ = _0921_ & _0122_;
  assign _0433_ = _0923_ & _0124_;
  assign _0436_ = _0925_ & _0126_;
  assign _0425_ = _0911_ & _0913_;
  assign _0428_ = _0915_ & _0917_;
  assign _0431_ = _0919_ & _0921_;
  assign _0434_ = _0938_ & _0923_;
  assign _0437_ = _0940_ & _0925_;
  assign _0745_ = _0423_ | _0424_;
  assign _0746_ = _0426_ | _0427_;
  assign _0747_ = _0429_ | _0430_;
  assign _0748_ = _0432_ | _0433_;
  assign _0749_ = _0435_ | _0436_;
  assign _0935_ = _0745_ | _0425_;
  assign _0005_ = _0746_ | _0428_;
  assign _0938_ = _0747_ | _0431_;
  assign _0940_ = _0748_ | _0434_;
  assign _0043_ = _0749_ | _0437_;
  assign _0102_ = ~ { _0979_, _0979_, _0979_, _0979_, _0979_, _0979_, _0979_, _0979_, _0979_, _0979_, _0979_, _0979_, _0979_, _0979_, _0979_, _0979_, _0979_, _0979_, _0979_, _0979_, _0979_, _0979_, _0979_, _0979_, _0979_, _0979_, _0979_, _0979_, _0979_, _0979_, _0979_, _0979_ };
  assign _0103_ = ~ { _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_ };
  assign _0104_ = ~ { _0983_, _0983_, _0983_, _0983_, _0983_, _0983_, _0983_, _0983_, _0983_, _0983_, _0983_, _0983_, _0983_, _0983_, _0983_, _0983_, _0983_, _0983_, _0983_, _0983_, _0983_, _0983_, _0983_, _0983_, _0983_, _0983_, _0983_, _0983_, _0983_, _0983_, _0983_, _0983_ };
  assign _0105_ = ~ { _0637_, _0637_, _0637_, _0637_, _0637_, _0637_, _0637_, _0637_, _0637_, _0637_, _0637_, _0637_, _0637_, _0637_, _0637_, _0637_, _0637_, _0637_, _0637_, _0637_, _0637_, _0637_, _0637_, _0637_, _0637_, _0637_, _0637_, _0637_, _0637_, _0637_, _0637_, _0637_ };
  assign _0106_ = ~ { _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_ };
  assign _0107_ = ~ { _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_ };
  assign _0108_ = ~ { _0639_, _0639_, _0639_, _0639_, _0639_, _0639_, _0639_, _0639_, _0639_, _0639_, _0639_, _0639_, _0639_, _0639_, _0639_, _0639_, _0639_, _0639_, _0639_, _0639_, _0639_, _0639_, _0639_, _0639_, _0639_, _0639_, _0639_, _0639_, _0639_, _0639_, _0639_, _0639_ };
  assign _0109_ = ~ id_fsm_q;
  assign _0110_ = ~ { rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel };
  assign _0111_ = ~ { _1021_, _1021_, _1021_, _1021_, _1021_, _1021_, _1021_, _1021_, _1021_, _1021_, _1021_, _1021_, _1021_, _1021_, _1021_, _1021_, _1021_, _1021_, _1021_, _1021_, _1021_, _1021_, _1021_, _1021_, _1021_, _1021_, _1021_, _1021_, _1021_, _1021_, _1021_, _1021_ };
  assign _0112_ = ~ { _1025_, _1025_, _1025_, _1025_, _1025_, _1025_, _1025_, _1025_, _1025_, _1025_, _1025_, _1025_, _1025_, _1025_, _1025_, _1025_, _1025_, _1025_, _1025_, _1025_, _1025_, _1025_, _1025_, _1025_, _1025_, _1025_, _1025_, _1025_, _1025_, _1025_, _1025_, _1025_ };
  assign _0113_ = ~ { _0641_, _0641_, _0641_, _0641_, _0641_, _0641_, _0641_, _0641_, _0641_, _0641_, _0641_, _0641_, _0641_, _0641_, _0641_, _0641_, _0641_, _0641_, _0641_, _0641_, _0641_, _0641_, _0641_, _0641_, _0641_, _0641_, _0641_, _0641_, _0641_, _0641_, _0641_, _0641_ };
  assign _0158_ = ~ { _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_ };
  assign _0160_ = ~ _0070_;
  assign _0162_ = ~ lsu_req_done_i;
  assign _0163_ = ~ alu_multicycle_dec;
  assign _0166_ = ~ jump_in_dec;
  assign _0164_ = ~ branch_in_dec;
  assign _0161_ = ~ multdiv_en_dec;
  assign _0165_ = ~ lsu_req_dec;
  assign _0167_ = ~ instr_executing_spec;
  assign _0168_ = ~ _0930_;
  assign _0172_ = ~ { lsu_addr_incr_req_i, lsu_addr_incr_req_i };
  assign _0173_ = ~ lsu_addr_incr_req_i;
  assign _0174_ = ~ { lsu_addr_incr_req_i, lsu_addr_incr_req_i, lsu_addr_incr_req_i };
  assign _0175_ = ~ { imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel };
  assign _0176_ = ~ { instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i };
  assign _0177_ = ~ { alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel };
  assign _0137_ = ~ data_ind_timing_i;
  assign _0178_ = ~ { _0081_, _0081_, _0081_, _0081_, _0081_, _0081_, _0081_, _0081_, _0081_, _0081_, _0081_, _0081_, _0081_, _0081_, _0081_, _0081_, _0081_, _0081_, _0081_, _0081_, _0081_, _0081_, _0081_, _0081_, _0081_, _0081_, _0081_, _0081_, _0081_, _0081_, _0081_, _0081_ };
  assign _0179_ = ~ { _0083_, _0083_, _0083_, _0083_, _0083_, _0083_, _0083_, _0083_, _0083_, _0083_, _0083_, _0083_, _0083_, _0083_, _0083_, _0083_, _0083_, _0083_, _0083_, _0083_, _0083_, _0083_, _0083_, _0083_, _0083_, _0083_, _0083_, _0083_, _0083_, _0083_, _0083_, _0083_ };
  assign _0180_ = ~ { lsu_we_o, lsu_we_o };
  assign _0181_ = ~ { lsu_req_dec, lsu_req_dec };
  assign _0702_ = { _0980_, _0980_, _0980_, _0980_, _0980_, _0980_, _0980_, _0980_, _0980_, _0980_, _0980_, _0980_, _0980_, _0980_, _0980_, _0980_, _0980_, _0980_, _0980_, _0980_, _0980_, _0980_, _0980_, _0980_, _0980_, _0980_, _0980_, _0980_, _0980_, _0980_, _0980_, _0980_ } | _0102_;
  assign _0705_ = { _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_ } | _0103_;
  assign _0708_ = { _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_ } | _0104_;
  assign _0711_ = { _0638_, _0638_, _0638_, _0638_, _0638_, _0638_, _0638_, _0638_, _0638_, _0638_, _0638_, _0638_, _0638_, _0638_, _0638_, _0638_, _0638_, _0638_, _0638_, _0638_, _0638_, _0638_, _0638_, _0638_, _0638_, _0638_, _0638_, _0638_, _0638_, _0638_, _0638_, _0638_ } | _0105_;
  assign _0714_ = { _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_ } | _0106_;
  assign _0717_ = { _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_ } | _0107_;
  assign _0720_ = { _0640_, _0640_, _0640_, _0640_, _0640_, _0640_, _0640_, _0640_, _0640_, _0640_, _0640_, _0640_, _0640_, _0640_, _0640_, _0640_, _0640_, _0640_, _0640_, _0640_, _0640_, _0640_, _0640_, _0640_, _0640_, _0640_, _0640_, _0640_, _0640_, _0640_, _0640_, _0640_ } | _0108_;
  assign _0723_ = id_fsm_q_t0 | _0109_;
  assign _0729_ = { rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0 } | _0110_;
  assign _0732_ = { _1022_, _1022_, _1022_, _1022_, _1022_, _1022_, _1022_, _1022_, _1022_, _1022_, _1022_, _1022_, _1022_, _1022_, _1022_, _1022_, _1022_, _1022_, _1022_, _1022_, _1022_, _1022_, _1022_, _1022_, _1022_, _1022_, _1022_, _1022_, _1022_, _1022_, _1022_, _1022_ } | _0111_;
  assign _0735_ = { _1026_, _1026_, _1026_, _1026_, _1026_, _1026_, _1026_, _1026_, _1026_, _1026_, _1026_, _1026_, _1026_, _1026_, _1026_, _1026_, _1026_, _1026_, _1026_, _1026_, _1026_, _1026_, _1026_, _1026_, _1026_, _1026_, _1026_, _1026_, _1026_, _1026_, _1026_, _1026_ } | _0112_;
  assign _0738_ = { _0642_, _0642_, _0642_, _0642_, _0642_, _0642_, _0642_, _0642_, _0642_, _0642_, _0642_, _0642_, _0642_, _0642_, _0642_, _0642_, _0642_, _0642_, _0642_, _0642_, _0642_, _0642_, _0642_, _0642_, _0642_, _0642_, _0642_, _0642_, _0642_, _0642_, _0642_, _0642_ } | _0113_;
  assign _0766_ = { _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_ } | _0158_;
  assign _0769_ = _0057_ | _0160_;
  assign _0774_ = alu_multicycle_dec_t0 | _0163_;
  assign _0782_ = jump_in_dec_t0 | _0166_;
  assign _0770_ = multdiv_en_dec_t0 | _0161_;
  assign _0779_ = lsu_req_dec_t0 | _0165_;
  assign _0775_ = branch_in_dec_t0 | _0164_;
  assign _0788_ = instr_executing_spec_t0 | _0167_;
  assign _0792_ = _0931_ | _0168_;
  assign _0795_ = { lsu_addr_incr_req_i_t0, lsu_addr_incr_req_i_t0 } | _0172_;
  assign _0798_ = lsu_addr_incr_req_i_t0 | _0173_;
  assign _0799_ = { lsu_addr_incr_req_i_t0, lsu_addr_incr_req_i_t0, lsu_addr_incr_req_i_t0 } | _0174_;
  assign _0802_ = { imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0 } | _0175_;
  assign _0805_ = { instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0 } | _0176_;
  assign _0808_ = { alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0 } | _0177_;
  assign _0813_ = { _0082_, _0082_, _0082_, _0082_, _0082_, _0082_, _0082_, _0082_, _0082_, _0082_, _0082_, _0082_, _0082_, _0082_, _0082_, _0082_, _0082_, _0082_, _0082_, _0082_, _0082_, _0082_, _0082_, _0082_, _0082_, _0082_, _0082_, _0082_, _0082_, _0082_, _0082_, _0082_ } | _0178_;
  assign _0816_ = { _0084_, _0084_, _0084_, _0084_, _0084_, _0084_, _0084_, _0084_, _0084_, _0084_, _0084_, _0084_, _0084_, _0084_, _0084_, _0084_, _0084_, _0084_, _0084_, _0084_, _0084_, _0084_, _0084_, _0084_, _0084_, _0084_, _0084_, _0084_, _0084_, _0084_, _0084_, _0084_ } | _0179_;
  assign _0819_ = { lsu_we_o_t0, lsu_we_o_t0 } | _0180_;
  assign _0822_ = { lsu_req_dec_t0, lsu_req_dec_t0 } | _0181_;
  assign _0703_ = { _0980_, _0980_, _0980_, _0980_, _0980_, _0980_, _0980_, _0980_, _0980_, _0980_, _0980_, _0980_, _0980_, _0980_, _0980_, _0980_, _0980_, _0980_, _0980_, _0980_, _0980_, _0980_, _0980_, _0980_, _0980_, _0980_, _0980_, _0980_, _0980_, _0980_, _0980_, _0980_ } | { _0979_, _0979_, _0979_, _0979_, _0979_, _0979_, _0979_, _0979_, _0979_, _0979_, _0979_, _0979_, _0979_, _0979_, _0979_, _0979_, _0979_, _0979_, _0979_, _0979_, _0979_, _0979_, _0979_, _0979_, _0979_, _0979_, _0979_, _0979_, _0979_, _0979_, _0979_, _0979_ };
  assign _0706_ = { _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_ } | { _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_ };
  assign _0709_ = { _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_ } | { _0983_, _0983_, _0983_, _0983_, _0983_, _0983_, _0983_, _0983_, _0983_, _0983_, _0983_, _0983_, _0983_, _0983_, _0983_, _0983_, _0983_, _0983_, _0983_, _0983_, _0983_, _0983_, _0983_, _0983_, _0983_, _0983_, _0983_, _0983_, _0983_, _0983_, _0983_, _0983_ };
  assign _0712_ = { _0638_, _0638_, _0638_, _0638_, _0638_, _0638_, _0638_, _0638_, _0638_, _0638_, _0638_, _0638_, _0638_, _0638_, _0638_, _0638_, _0638_, _0638_, _0638_, _0638_, _0638_, _0638_, _0638_, _0638_, _0638_, _0638_, _0638_, _0638_, _0638_, _0638_, _0638_, _0638_ } | { _0637_, _0637_, _0637_, _0637_, _0637_, _0637_, _0637_, _0637_, _0637_, _0637_, _0637_, _0637_, _0637_, _0637_, _0637_, _0637_, _0637_, _0637_, _0637_, _0637_, _0637_, _0637_, _0637_, _0637_, _0637_, _0637_, _0637_, _0637_, _0637_, _0637_, _0637_, _0637_ };
  assign _0715_ = { _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_ } | { _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_ };
  assign _0718_ = { _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_ } | { _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_ };
  assign _0721_ = { _0640_, _0640_, _0640_, _0640_, _0640_, _0640_, _0640_, _0640_, _0640_, _0640_, _0640_, _0640_, _0640_, _0640_, _0640_, _0640_, _0640_, _0640_, _0640_, _0640_, _0640_, _0640_, _0640_, _0640_, _0640_, _0640_, _0640_, _0640_, _0640_, _0640_, _0640_, _0640_ } | { _0639_, _0639_, _0639_, _0639_, _0639_, _0639_, _0639_, _0639_, _0639_, _0639_, _0639_, _0639_, _0639_, _0639_, _0639_, _0639_, _0639_, _0639_, _0639_, _0639_, _0639_, _0639_, _0639_, _0639_, _0639_, _0639_, _0639_, _0639_, _0639_, _0639_, _0639_, _0639_ };
  assign _0724_ = id_fsm_q_t0 | id_fsm_q;
  assign _0730_ = { rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0 } | { rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel };
  assign _0733_ = { _1022_, _1022_, _1022_, _1022_, _1022_, _1022_, _1022_, _1022_, _1022_, _1022_, _1022_, _1022_, _1022_, _1022_, _1022_, _1022_, _1022_, _1022_, _1022_, _1022_, _1022_, _1022_, _1022_, _1022_, _1022_, _1022_, _1022_, _1022_, _1022_, _1022_, _1022_, _1022_ } | { _1021_, _1021_, _1021_, _1021_, _1021_, _1021_, _1021_, _1021_, _1021_, _1021_, _1021_, _1021_, _1021_, _1021_, _1021_, _1021_, _1021_, _1021_, _1021_, _1021_, _1021_, _1021_, _1021_, _1021_, _1021_, _1021_, _1021_, _1021_, _1021_, _1021_, _1021_, _1021_ };
  assign _0736_ = { _1026_, _1026_, _1026_, _1026_, _1026_, _1026_, _1026_, _1026_, _1026_, _1026_, _1026_, _1026_, _1026_, _1026_, _1026_, _1026_, _1026_, _1026_, _1026_, _1026_, _1026_, _1026_, _1026_, _1026_, _1026_, _1026_, _1026_, _1026_, _1026_, _1026_, _1026_, _1026_ } | { _1025_, _1025_, _1025_, _1025_, _1025_, _1025_, _1025_, _1025_, _1025_, _1025_, _1025_, _1025_, _1025_, _1025_, _1025_, _1025_, _1025_, _1025_, _1025_, _1025_, _1025_, _1025_, _1025_, _1025_, _1025_, _1025_, _1025_, _1025_, _1025_, _1025_, _1025_, _1025_ };
  assign _0739_ = { _0642_, _0642_, _0642_, _0642_, _0642_, _0642_, _0642_, _0642_, _0642_, _0642_, _0642_, _0642_, _0642_, _0642_, _0642_, _0642_, _0642_, _0642_, _0642_, _0642_, _0642_, _0642_, _0642_, _0642_, _0642_, _0642_, _0642_, _0642_, _0642_, _0642_, _0642_, _0642_ } | { _0641_, _0641_, _0641_, _0641_, _0641_, _0641_, _0641_, _0641_, _0641_, _0641_, _0641_, _0641_, _0641_, _0641_, _0641_, _0641_, _0641_, _0641_, _0641_, _0641_, _0641_, _0641_, _0641_, _0641_, _0641_, _0641_, _0641_, _0641_, _0641_, _0641_, _0641_, _0641_ };
  assign _0767_ = { _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_ } | { _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_ };
  assign _0773_ = ex_valid_i_t0 | ex_valid_i;
  assign _0783_ = jump_in_dec_t0 | jump_in_dec;
  assign _0776_ = branch_in_dec_t0 | branch_in_dec;
  assign _0771_ = multdiv_en_dec_t0 | multdiv_en_dec;
  assign _0780_ = lsu_req_dec_t0 | lsu_req_dec;
  assign _0789_ = instr_executing_spec_t0 | instr_executing_spec;
  assign _0791_ = _0933_ | _0932_;
  assign _0793_ = _0931_ | _0930_;
  assign _0796_ = { lsu_addr_incr_req_i_t0, lsu_addr_incr_req_i_t0 } | { lsu_addr_incr_req_i, lsu_addr_incr_req_i };
  assign _0800_ = { lsu_addr_incr_req_i_t0, lsu_addr_incr_req_i_t0, lsu_addr_incr_req_i_t0 } | { lsu_addr_incr_req_i, lsu_addr_incr_req_i, lsu_addr_incr_req_i };
  assign _0803_ = { imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0 } | { imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel };
  assign _0806_ = { instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0 } | { instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i };
  assign _0809_ = { alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0 } | { alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel };
  assign _0811_ = instr_executing_t0 | instr_executing;
  assign _0814_ = { _0082_, _0082_, _0082_, _0082_, _0082_, _0082_, _0082_, _0082_, _0082_, _0082_, _0082_, _0082_, _0082_, _0082_, _0082_, _0082_, _0082_, _0082_, _0082_, _0082_, _0082_, _0082_, _0082_, _0082_, _0082_, _0082_, _0082_, _0082_, _0082_, _0082_, _0082_, _0082_ } | { _0081_, _0081_, _0081_, _0081_, _0081_, _0081_, _0081_, _0081_, _0081_, _0081_, _0081_, _0081_, _0081_, _0081_, _0081_, _0081_, _0081_, _0081_, _0081_, _0081_, _0081_, _0081_, _0081_, _0081_, _0081_, _0081_, _0081_, _0081_, _0081_, _0081_, _0081_, _0081_ };
  assign _0817_ = { _0084_, _0084_, _0084_, _0084_, _0084_, _0084_, _0084_, _0084_, _0084_, _0084_, _0084_, _0084_, _0084_, _0084_, _0084_, _0084_, _0084_, _0084_, _0084_, _0084_, _0084_, _0084_, _0084_, _0084_, _0084_, _0084_, _0084_, _0084_, _0084_, _0084_, _0084_, _0084_ } | { _0083_, _0083_, _0083_, _0083_, _0083_, _0083_, _0083_, _0083_, _0083_, _0083_, _0083_, _0083_, _0083_, _0083_, _0083_, _0083_, _0083_, _0083_, _0083_, _0083_, _0083_, _0083_, _0083_, _0083_, _0083_, _0083_, _0083_, _0083_, _0083_, _0083_, _0083_, _0083_ };
  assign _0820_ = { lsu_we_o_t0, lsu_we_o_t0 } | { lsu_we_o, lsu_we_o };
  assign _0823_ = { lsu_req_dec_t0, lsu_req_dec_t0 } | { lsu_req_dec, lsu_req_dec };
  assign _0346_ = imm_u_type_t0 & _0702_;
  assign _0349_ = 32'd0 & _0705_;
  assign _0352_ = _0899_ & _0708_;
  assign _0355_ = _0901_ & _0711_;
  assign _0358_ = imm_b_type_t0 & _0714_;
  assign _0361_ = _1032_ & _0717_;
  assign _0364_ = _0905_ & _0720_;
  assign _0367_ = _0029_ & _0723_;
  assign _0370_ = _0037_ & _0723_;
  assign _0372_ = _0035_ & _0723_;
  assign _0377_ = _0039_ & _0723_;
  assign _0380_ = _0041_ & _0723_;
  assign _0383_ = _0031_ & _0723_;
  assign _0385_ = _0023_ & _0723_;
  assign _0387_ = _0025_ & _0723_;
  assign _0389_ = _0033_ & _0723_;
  assign _0391_ = result_ex_i_t0 & _0729_;
  assign _0394_ = pc_id_i_t0 & _0732_;
  assign _0397_ = multdiv_operand_a_ex_o_t0 & _0735_;
  assign _0400_ = _0909_ & _0738_;
  assign _0493_ = pc_id_i_t0 & _0766_;
  assign _0497_ = jump_in_dec_t0 & _0769_;
  assign _0499_ = branch_in_dec_t0 & _0769_;
  assign _0501_ = multdiv_en_dec_t0 & _0769_;
  assign _0503_ = rf_we_dec_t0 & _0770_;
  assign _0510_ = _0997_ & _0770_;
  assign _0513_ = _0999_ & _0779_;
  assign _0516_ = alu_multicycle_dec_t0 & _0782_;
  assign _0507_ = _0995_ & _0775_;
  assign _0519_ = _1000_ & _0770_;
  assign _0521_ = _1001_ & _0779_;
  assign _0523_ = rf_we_dec_t0 & _0774_;
  assign _0525_ = _1003_ & _0782_;
  assign _0528_ = _1005_ & _0775_;
  assign _0531_ = _1007_ & _0770_;
  assign _0534_ = _1009_ & _0779_;
  assign _0538_ = _1010_ & _0770_;
  assign _0540_ = _1011_ & _0779_;
  assign _0543_ = _1012_ & _0779_;
  assign _0547_ = _1013_ & _0775_;
  assign _0549_ = _1014_ & _0770_;
  assign _0551_ = _1015_ & _0779_;
  assign _0555_ = _1016_ & _0770_;
  assign _0557_ = _1017_ & _0779_;
  assign _0561_ = _1018_ & _0770_;
  assign _0563_ = _1019_ & _0779_;
  assign _0565_ = branch_in_dec_t0 & _0770_;
  assign _0567_ = _1020_ & _0779_;
  assign _0571_ = rf_we_dec_t0 & _0788_;
  assign _0590_ = _0027_ & _0792_;
  assign _0599_ = alu_op_a_mux_sel_dec_t0 & _0795_;
  assign _0602_ = alu_op_b_mux_sel_dec_t0 & _0798_;
  assign _0604_ = imm_b_mux_sel_dec_t0 & _0799_;
  assign _0607_ = zimm_rs1_type_t0 & _0802_;
  assign _0610_ = 32'd0 & _0805_;
  assign _0613_ = lsu_wdata_o_t0 & _0808_;
  assign _0622_ = ex_valid_i_t0 & _0779_;
  assign _0625_ = rf_rdata_a_i_t0 & _0813_;
  assign _0628_ = rf_rdata_b_i_t0 & _0816_;
  assign _0631_ = 2'h0 & _0819_;
  assign _0634_ = 2'h0 & _0822_;
  assign _0347_ = _1032_ & _0703_;
  assign _0350_ = imm_i_type_t0 & _0706_;
  assign _0353_ = imm_s_type_t0 & _0709_;
  assign _0356_ = _0897_ & _0712_;
  assign _0359_ = imm_j_type_t0 & _0715_;
  assign _0362_ = imm_i_type_t0 & _0718_;
  assign _0365_ = _0903_ & _0721_;
  assign _0368_ = _0057_ & _0724_;
  assign _0373_ = _0053_ & _0724_;
  assign _0375_ = _0050_ & _0724_;
  assign _0378_ = _0048_ & _0724_;
  assign _0381_ = _0055_ & _0724_;
  assign _0392_ = csr_rdata_i_t0 & _0730_;
  assign _0395_ = imm_a_t0 & _0733_;
  assign _0398_ = lsu_addr_last_i_t0 & _0736_;
  assign _0401_ = _0907_ & _0739_;
  assign _0494_ = multdiv_operand_a_ex_o_t0 & _0767_;
  assign _0504_ = _0069_ & _0771_;
  assign _0506_ = rf_we_dec_t0 & _0773_;
  assign _0514_ = lsu_req_done_i_t0 & _0780_;
  assign _0526_ = rf_we_dec_t0 & _0783_;
  assign _0529_ = rf_we_dec_t0 & _0776_;
  assign _0532_ = _0046_ & _0771_;
  assign _0535_ = rf_we_dec_t0 & _0780_;
  assign _0508_ = data_ind_timing_i_t0 & _0776_;
  assign _0511_ = ex_valid_i_t0 & _0771_;
  assign _0545_ = jump_set_dec_t0 & _0783_;
  assign _0553_ = _0960_ & _0776_;
  assign _0559_ = branch_decision_i_t0 & _0776_;
  assign _0569_ = _0015_ & _0789_;
  assign _0572_ = _0013_ & _0789_;
  assign _0574_ = _0019_ & _0789_;
  assign _0576_ = _0017_ & _0789_;
  assign _0578_ = _0021_ & _0789_;
  assign _0580_ = _0009_ & _0789_;
  assign _0582_ = _0001_ & _0789_;
  assign _0584_ = _0003_ & _0789_;
  assign _0586_ = _0011_ & _0789_;
  assign _0588_ = _0043_ & _0791_;
  assign _0591_ = _0005_ & _0793_;
  assign _0600_ = 2'h0 & _0796_;
  assign _0605_ = 3'h0 & _0800_;
  assign _0608_ = 32'd0 & _0803_;
  assign _0611_ = 32'd0 & _0806_;
  assign _0614_ = imm_b_t0 & _0809_;
  assign _0616_ = _0065_ & _0811_;
  assign _0618_ = mult_en_dec_t0 & _0811_;
  assign _0620_ = div_en_dec_t0 & _0811_;
  assign _0623_ = stall_mem_t0 & _0780_;
  assign _0626_ = rf_wdata_fwd_wb_i_t0 & _0814_;
  assign _0629_ = rf_wdata_fwd_wb_i_t0 & _0817_;
  assign _0632_ = 2'h0 & _0820_;
  assign _0635_ = _1035_ & _0823_;
  assign _0704_ = _0346_ | _0347_;
  assign _0707_ = _0349_ | _0350_;
  assign _0710_ = _0352_ | _0353_;
  assign _0713_ = _0355_ | _0356_;
  assign _0716_ = _0358_ | _0359_;
  assign _0719_ = _0361_ | _0362_;
  assign _0722_ = _0364_ | _0365_;
  assign _0725_ = _0367_ | _0368_;
  assign _0726_ = _0372_ | _0373_;
  assign _0727_ = _0377_ | _0378_;
  assign _0728_ = _0380_ | _0381_;
  assign _0731_ = _0391_ | _0392_;
  assign _0734_ = _0394_ | _0395_;
  assign _0737_ = _0397_ | _0398_;
  assign _0740_ = _0400_ | _0401_;
  assign _0768_ = _0493_ | _0494_;
  assign _0772_ = _0503_ | _0504_;
  assign _0777_ = _0507_ | _0508_;
  assign _0778_ = _0510_ | _0511_;
  assign _0781_ = _0513_ | _0514_;
  assign _0784_ = _0525_ | _0526_;
  assign _0785_ = _0528_ | _0529_;
  assign _0786_ = _0531_ | _0532_;
  assign _0787_ = _0534_ | _0535_;
  assign _0790_ = _0571_ | _0572_;
  assign _0794_ = _0590_ | _0591_;
  assign _0797_ = _0599_ | _0600_;
  assign _0801_ = _0604_ | _0605_;
  assign _0804_ = _0607_ | _0608_;
  assign _0807_ = _0610_ | _0611_;
  assign _0810_ = _0613_ | _0614_;
  assign _0812_ = _0622_ | _0623_;
  assign _0815_ = _0625_ | _0626_;
  assign _0818_ = _0628_ | _0629_;
  assign _0821_ = _0631_ | _0632_;
  assign _0824_ = _0634_ | _0635_;
  assign _0828_ = imm_u_type ^ _1031_;
  assign _0829_ = 32'd4 ^ imm_i_type;
  assign _0830_ = _0898_ ^ imm_s_type;
  assign _0831_ = _0900_ ^ _0896_;
  assign _0832_ = imm_b_type ^ imm_j_type;
  assign _0833_ = _1031_ ^ imm_i_type;
  assign _0834_ = _0904_ ^ _0902_;
  assign _0835_ = _0028_ ^ _0056_;
  assign _0836_ = _0034_ ^ _0052_;
  assign _0837_ = _0038_ ^ _0047_;
  assign _0838_ = _0040_ ^ _0054_;
  assign _0839_ = result_ex_i ^ csr_rdata_i;
  assign _0840_ = pc_id_i ^ imm_a;
  assign _0841_ = multdiv_operand_a_ex_o ^ lsu_addr_last_i;
  assign _0842_ = _0908_ ^ _0906_;
  assign _0843_ = pc_id_i ^ multdiv_operand_a_ex_o;
  assign _0844_ = rf_we_dec ^ _0068_;
  assign _0845_ = _0849_ ^ _1033_;
  assign _0846_ = _0996_ ^ _0051_;
  assign _0847_ = _0998_ ^ _0044_;
  assign _0852_ = _1002_ ^ rf_we_dec;
  assign _0853_ = _1004_ ^ rf_we_dec;
  assign _0854_ = _1006_ ^ _0045_;
  assign _0855_ = _1008_ ^ rf_we_dec;
  assign _0869_ = rf_we_dec ^ _0012_;
  assign _0870_ = _0026_ ^ _0004_;
  assign _0871_ = alu_op_a_mux_sel_dec ^ 2'h1;
  assign _0872_ = imm_b_mux_sel_dec ^ 3'h6;
  assign _0873_ = lsu_wdata_o ^ imm_b;
  assign _0874_ = ex_valid_i ^ _0139_;
  assign _0875_ = rf_rdata_a_i ^ rf_wdata_fwd_wb_i;
  assign _0876_ = rf_rdata_b_i ^ rf_wdata_fwd_wb_i;
  assign _0877_ = 2'h2 ^ _1034_;
  assign _0348_ = { _0980_, _0980_, _0980_, _0980_, _0980_, _0980_, _0980_, _0980_, _0980_, _0980_, _0980_, _0980_, _0980_, _0980_, _0980_, _0980_, _0980_, _0980_, _0980_, _0980_, _0980_, _0980_, _0980_, _0980_, _0980_, _0980_, _0980_, _0980_, _0980_, _0980_, _0980_, _0980_ } & _0828_;
  assign _0351_ = { _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_ } & _0829_;
  assign _0354_ = { _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_ } & _0830_;
  assign _0357_ = { _0638_, _0638_, _0638_, _0638_, _0638_, _0638_, _0638_, _0638_, _0638_, _0638_, _0638_, _0638_, _0638_, _0638_, _0638_, _0638_, _0638_, _0638_, _0638_, _0638_, _0638_, _0638_, _0638_, _0638_, _0638_, _0638_, _0638_, _0638_, _0638_, _0638_, _0638_, _0638_ } & _0831_;
  assign _0360_ = { _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_ } & _0832_;
  assign _0363_ = { _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_ } & _0833_;
  assign _0366_ = { _0640_, _0640_, _0640_, _0640_, _0640_, _0640_, _0640_, _0640_, _0640_, _0640_, _0640_, _0640_, _0640_, _0640_, _0640_, _0640_, _0640_, _0640_, _0640_, _0640_, _0640_, _0640_, _0640_, _0640_, _0640_, _0640_, _0640_, _0640_, _0640_, _0640_, _0640_, _0640_ } & _0834_;
  assign _0369_ = id_fsm_q_t0 & _0835_;
  assign _0371_ = id_fsm_q_t0 & _0036_;
  assign _0374_ = id_fsm_q_t0 & _0836_;
  assign _0376_ = id_fsm_q_t0 & _0049_;
  assign _0379_ = id_fsm_q_t0 & _0837_;
  assign _0382_ = id_fsm_q_t0 & _0838_;
  assign _0384_ = id_fsm_q_t0 & _0030_;
  assign _0386_ = id_fsm_q_t0 & _0022_;
  assign _0388_ = id_fsm_q_t0 & _0024_;
  assign _0390_ = id_fsm_q_t0 & _0032_;
  assign _0393_ = { rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0 } & _0839_;
  assign _0396_ = { _1022_, _1022_, _1022_, _1022_, _1022_, _1022_, _1022_, _1022_, _1022_, _1022_, _1022_, _1022_, _1022_, _1022_, _1022_, _1022_, _1022_, _1022_, _1022_, _1022_, _1022_, _1022_, _1022_, _1022_, _1022_, _1022_, _1022_, _1022_, _1022_, _1022_, _1022_, _1022_ } & _0840_;
  assign _0399_ = { _1026_, _1026_, _1026_, _1026_, _1026_, _1026_, _1026_, _1026_, _1026_, _1026_, _1026_, _1026_, _1026_, _1026_, _1026_, _1026_, _1026_, _1026_, _1026_, _1026_, _1026_, _1026_, _1026_, _1026_, _1026_, _1026_, _1026_, _1026_, _1026_, _1026_, _1026_, _1026_ } & _0841_;
  assign _0402_ = { _0642_, _0642_, _0642_, _0642_, _0642_, _0642_, _0642_, _0642_, _0642_, _0642_, _0642_, _0642_, _0642_, _0642_, _0642_, _0642_, _0642_, _0642_, _0642_, _0642_, _0642_, _0642_, _0642_, _0642_, _0642_, _0642_, _0642_, _0642_, _0642_, _0642_, _0642_, _0642_ } & _0842_;
  assign _0495_ = { _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_ } & _0843_;
  assign _0498_ = _0057_ & jump_in_dec;
  assign _0500_ = _0057_ & branch_in_dec;
  assign _0502_ = _0057_ & multdiv_en_dec;
  assign _0505_ = multdiv_en_dec_t0 & _0844_;
  assign _0241_ = ex_valid_i_t0 & rf_we_dec;
  assign _0509_ = branch_in_dec_t0 & _0845_;
  assign _0512_ = multdiv_en_dec_t0 & _0846_;
  assign _0515_ = lsu_req_dec_t0 & _0847_;
  assign _0517_ = jump_in_dec_t0 & _0848_;
  assign _0518_ = branch_in_dec_t0 & _0849_;
  assign _0520_ = multdiv_en_dec_t0 & _0850_;
  assign _0522_ = lsu_req_dec_t0 & _0851_;
  assign _0524_ = alu_multicycle_dec_t0 & rf_we_dec;
  assign _0527_ = jump_in_dec_t0 & _0852_;
  assign _0530_ = branch_in_dec_t0 & _0853_;
  assign _0533_ = multdiv_en_dec_t0 & _0854_;
  assign _0536_ = lsu_req_dec_t0 & _0855_;
  assign _0537_ = branch_in_dec_t0 & data_ind_timing_i;
  assign _0539_ = multdiv_en_dec_t0 & _0856_;
  assign _0541_ = lsu_req_dec_t0 & _0857_;
  assign _0542_ = multdiv_en_dec_t0 & _0051_;
  assign _0544_ = lsu_req_dec_t0 & _0858_;
  assign _0546_ = jump_in_dec_t0 & jump_set_dec;
  assign _0548_ = branch_in_dec_t0 & _0859_;
  assign _0550_ = multdiv_en_dec_t0 & _0860_;
  assign _0552_ = lsu_req_dec_t0 & _0861_;
  assign _0554_ = branch_in_dec_t0 & _0862_;
  assign _0556_ = multdiv_en_dec_t0 & _0863_;
  assign _0558_ = lsu_req_dec_t0 & _0864_;
  assign _0560_ = branch_in_dec_t0 & branch_decision_i;
  assign _0562_ = multdiv_en_dec_t0 & _0865_;
  assign _0564_ = lsu_req_dec_t0 & _0866_;
  assign _0566_ = multdiv_en_dec_t0 & _0867_;
  assign _0568_ = lsu_req_dec_t0 & _0868_;
  assign _0570_ = instr_executing_spec_t0 & _0014_;
  assign _0573_ = instr_executing_spec_t0 & _0869_;
  assign _0575_ = instr_executing_spec_t0 & _0018_;
  assign _0577_ = instr_executing_spec_t0 & _0016_;
  assign _0579_ = instr_executing_spec_t0 & _0020_;
  assign _0581_ = instr_executing_spec_t0 & _0008_;
  assign _0583_ = instr_executing_spec_t0 & _0000_;
  assign _0585_ = instr_executing_spec_t0 & _0002_;
  assign _0587_ = instr_executing_spec_t0 & _0010_;
  assign _0589_ = _0933_ & _0042_;
  assign _0592_ = _0931_ & _0870_;
  assign _0601_ = { lsu_addr_incr_req_i_t0, lsu_addr_incr_req_i_t0 } & _0871_;
  assign _0603_ = lsu_addr_incr_req_i_t0 & _0182_;
  assign _0606_ = { lsu_addr_incr_req_i_t0, lsu_addr_incr_req_i_t0, lsu_addr_incr_req_i_t0 } & _0872_;
  assign _0609_ = { imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0 } & zimm_rs1_type;
  assign _0612_ = { instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0 } & 32'd6;
  assign _0615_ = { alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0 } & _0873_;
  assign _0617_ = instr_executing_t0 & _0064_;
  assign _0619_ = instr_executing_t0 & mult_en_dec;
  assign _0621_ = instr_executing_t0 & div_en_dec;
  assign _0624_ = lsu_req_dec_t0 & _0874_;
  assign _0627_ = { _0082_, _0082_, _0082_, _0082_, _0082_, _0082_, _0082_, _0082_, _0082_, _0082_, _0082_, _0082_, _0082_, _0082_, _0082_, _0082_, _0082_, _0082_, _0082_, _0082_, _0082_, _0082_, _0082_, _0082_, _0082_, _0082_, _0082_, _0082_, _0082_, _0082_, _0082_, _0082_ } & _0875_;
  assign _0630_ = { _0084_, _0084_, _0084_, _0084_, _0084_, _0084_, _0084_, _0084_, _0084_, _0084_, _0084_, _0084_, _0084_, _0084_, _0084_, _0084_, _0084_, _0084_, _0084_, _0084_, _0084_, _0084_, _0084_, _0084_, _0084_, _0084_, _0084_, _0084_, _0084_, _0084_, _0084_, _0084_ } & _0876_;
  assign _0633_ = { lsu_we_o_t0, lsu_we_o_t0 } & 2'h1;
  assign _0636_ = { lsu_req_dec_t0, lsu_req_dec_t0 } & _0877_;
  assign _0897_ = _0348_ | _0704_;
  assign _0899_ = _0351_ | _0707_;
  assign _0901_ = _0354_ | _0710_;
  assign imm_b_t0 = _0357_ | _0713_;
  assign _0903_ = _0360_ | _0716_;
  assign _0905_ = _0363_ | _0719_;
  assign bt_b_operand_o_t0 = _0366_ | _0722_;
  assign _0007_ = _0369_ | _0725_;
  assign _0015_ = _0371_ | _0370_;
  assign _0013_ = _0374_ | _0726_;
  assign _0019_ = _0376_ | _0375_;
  assign _0017_ = _0379_ | _0727_;
  assign _0021_ = _0382_ | _0728_;
  assign _0009_ = _0384_ | _0383_;
  assign _0001_ = _0386_ | _0385_;
  assign _0003_ = _0388_ | _0387_;
  assign _0011_ = _0390_ | _0389_;
  assign rf_wdata_id_o_t0 = _0393_ | _0731_;
  assign _0907_ = _0396_ | _0734_;
  assign _0909_ = _0399_ | _0737_;
  assign alu_operand_a_ex_o_t0 = _0402_ | _0740_;
  assign bt_a_operand_o_t0 = _0495_ | _0768_;
  assign _0050_ = _0498_ | _0497_;
  assign _0048_ = _0500_ | _0499_;
  assign _0055_ = _0502_ | _0501_;
  assign _0053_ = _0505_ | _0772_;
  assign _0046_ = _0241_ | _0506_;
  assign _0997_ = _0509_ | _0777_;
  assign _0999_ = _0512_ | _0778_;
  assign _0029_ = _0515_ | _0781_;
  assign _0995_ = _0517_ | _0516_;
  assign _1000_ = _0518_ | _0507_;
  assign _1001_ = _0520_ | _0519_;
  assign _0037_ = _0522_ | _0521_;
  assign _1003_ = _0524_ | _0523_;
  assign _1005_ = _0527_ | _0784_;
  assign _1007_ = _0530_ | _0785_;
  assign _1009_ = _0533_ | _0786_;
  assign _0035_ = _0536_ | _0787_;
  assign _1010_ = _0537_ | _0508_;
  assign _1011_ = _0539_ | _0538_;
  assign _0039_ = _0541_ | _0540_;
  assign _1012_ = _0542_ | _0511_;
  assign _0041_ = _0544_ | _0543_;
  assign _1013_ = _0546_ | _0545_;
  assign _1014_ = _0548_ | _0547_;
  assign _1015_ = _0550_ | _0549_;
  assign _0031_ = _0552_ | _0551_;
  assign _1016_ = _0554_ | _0553_;
  assign _1017_ = _0556_ | _0555_;
  assign _0023_ = _0558_ | _0557_;
  assign _1018_ = _0560_ | _0559_;
  assign _1019_ = _0562_ | _0561_;
  assign _0025_ = _0564_ | _0563_;
  assign _1020_ = _0566_ | _0565_;
  assign _0033_ = _0568_ | _0567_;
  assign stall_alu_t0 = _0570_ | _0569_;
  assign rf_we_raw_t0 = _0573_ | _0790_;
  assign stall_jump_t0 = _0575_ | _0574_;
  assign stall_branch_t0 = _0577_ | _0576_;
  assign stall_multdiv_t0 = _0579_ | _0578_;
  assign jump_set_raw_t0 = _0581_ | _0580_;
  assign branch_set_raw_t0 = _0583_ | _0582_;
  assign branch_set_raw_spec_t0 = _0585_ | _0584_;
  assign perf_branch_o_t0 = _0587_ | _0586_;
  assign _0027_ = _0589_ | _0588_;
  assign csr_pipe_flush_t0 = _0592_ | _0794_;
  assign alu_op_a_mux_sel_t0 = _0601_ | _0797_;
  assign alu_op_b_mux_sel_t0 = _0603_ | _0602_;
  assign imm_b_mux_sel_t0 = _0606_ | _0801_;
  assign imm_a_t0 = _0609_ | _0804_;
  assign _1032_ = _0612_ | _0807_;
  assign alu_operand_b_ex_o_t0 = _0615_ | _0810_;
  assign lsu_req_o_t0 = _0617_ | _0616_;
  assign mult_en_ex_o_t0 = _0619_ | _0618_;
  assign div_en_ex_o_t0 = _0621_ | _0620_;
  assign multicycle_done_t0 = _0624_ | _0812_;
  assign multdiv_operand_a_ex_o_t0 = _0627_ | _0815_;
  assign lsu_wdata_o_t0 = _0630_ | _0818_;
  assign _1035_ = _0633_ | _0821_;
  assign instr_type_wb_o_t0 = _0636_ | _0824_;
  assign _0091_ = & { instr_executing, instr_executing_spec };
  assign _0182_ = ~ alu_op_b_mux_sel_dec;
  assign _0096_ = ~ _0981_;
  assign _0098_ = ~ _0989_;
  assign _0100_ = ~ _1023_;
  assign _0128_ = ~ illegal_insn_dec;
  assign _0130_ = ~ mult_en_dec;
  assign _0132_ = ~ branch_set_raw;
  assign _0134_ = ~ _0956_;
  assign _0136_ = ~ branch_decision_i;
  assign _0140_ = ~ _0961_;
  assign _0142_ = ~ _0963_;
  assign _0144_ = ~ _0965_;
  assign _0146_ = ~ _0967_;
  assign _0148_ = ~ outstanding_load_wb_i;
  assign _0150_ = ~ instr_fetch_err_i;
  assign _0152_ = ~ _0971_;
  assign _0154_ = ~ \gen_stall_mem.rf_rd_a_hz ;
  assign data_req_allowed = ~ \gen_stall_mem.outstanding_memory_access ;
  assign _0097_ = ~ _0979_;
  assign _0099_ = ~ _0987_;
  assign _0101_ = ~ _1021_;
  assign _0129_ = ~ illegal_csr_insn_i;
  assign _0131_ = ~ div_en_dec;
  assign _0133_ = ~ jump_set_raw;
  assign _0135_ = ~ branch_jump_set_done_q;
  assign _0139_ = ~ stall_mem;
  assign _0141_ = ~ stall_multdiv;
  assign _0143_ = ~ stall_jump;
  assign _0145_ = ~ stall_branch;
  assign _0147_ = ~ stall_alu;
  assign _0149_ = ~ outstanding_store_wb_i;
  assign _0151_ = ~ wb_exception;
  assign _0153_ = ~ _0079_;
  assign _0155_ = ~ \gen_stall_mem.rf_rd_b_hz ;
  assign _0138_ = ~ stall_ld_hz;
  assign _0337_ = _0982_ & _0097_;
  assign _0340_ = _0990_ & _0099_;
  assign _0343_ = _1024_ & _0101_;
  assign _0438_ = illegal_insn_dec_t0 & _0129_;
  assign _0441_ = mult_en_dec_t0 & _0131_;
  assign _0444_ = branch_set_raw_t0 & _0133_;
  assign _0447_ = _0957_ & _0135_;
  assign _0450_ = branch_decision_i_t0 & _0137_;
  assign _0453_ = stall_ld_hz_t0 & _0139_;
  assign _0456_ = _0962_ & _0141_;
  assign _0459_ = _0964_ & _0143_;
  assign _0462_ = _0966_ & _0145_;
  assign _0465_ = _0968_ & _0147_;
  assign _0468_ = outstanding_load_wb_i_t0 & _0149_;
  assign _0471_ = instr_fetch_err_i_t0 & _0151_;
  assign _0474_ = _0972_ & controller_run;
  assign _0477_ = data_req_allowed_t0 & _0153_;
  assign _0480_ = \gen_stall_mem.rf_rd_a_hz_t0  & _0155_;
  assign _0483_ = data_req_allowed_t0 & _0138_;
  assign _0338_ = _0980_ & _0096_;
  assign _0341_ = _0988_ & _0098_;
  assign _0344_ = _1022_ & _0100_;
  assign _0439_ = illegal_csr_insn_i_t0 & _0128_;
  assign _0442_ = div_en_dec_t0 & _0130_;
  assign _0445_ = jump_set_raw_t0 & _0132_;
  assign _0448_ = branch_jump_set_done_q_t0 & _0134_;
  assign _0451_ = data_ind_timing_i_t0 & _0136_;
  assign _0454_ = stall_mem_t0 & _0138_;
  assign _0457_ = stall_multdiv_t0 & _0140_;
  assign _0460_ = stall_jump_t0 & _0142_;
  assign _0463_ = stall_branch_t0 & _0144_;
  assign _0466_ = stall_alu_t0 & _0146_;
  assign _0469_ = outstanding_store_wb_i_t0 & _0148_;
  assign _0472_ = wb_exception_t0 & _0150_;
  assign _0475_ = controller_run_t0 & _0152_;
  assign _0478_ = _0080_ & data_req_allowed;
  assign _0481_ = \gen_stall_mem.rf_rd_b_hz_t0  & _0154_;
  assign _0484_ = stall_ld_hz_t0 & data_req_allowed;
  assign _0339_ = _0982_ & _0980_;
  assign _0342_ = _0990_ & _0988_;
  assign _0345_ = _1024_ & _1022_;
  assign _0440_ = illegal_insn_dec_t0 & illegal_csr_insn_i_t0;
  assign _0443_ = mult_en_dec_t0 & div_en_dec_t0;
  assign _0446_ = branch_set_raw_t0 & jump_set_raw_t0;
  assign _0449_ = _0957_ & branch_jump_set_done_q_t0;
  assign _0452_ = branch_decision_i_t0 & data_ind_timing_i_t0;
  assign _0455_ = stall_ld_hz_t0 & stall_mem_t0;
  assign _0458_ = _0962_ & stall_multdiv_t0;
  assign _0461_ = _0964_ & stall_jump_t0;
  assign _0464_ = _0966_ & stall_branch_t0;
  assign _0467_ = _0968_ & stall_alu_t0;
  assign _0470_ = outstanding_load_wb_i_t0 & outstanding_store_wb_i_t0;
  assign _0473_ = instr_fetch_err_i_t0 & wb_exception_t0;
  assign _0476_ = _0972_ & controller_run_t0;
  assign _0479_ = data_req_allowed_t0 & _0080_;
  assign _0482_ = \gen_stall_mem.rf_rd_a_hz_t0  & \gen_stall_mem.rf_rd_b_hz_t0 ;
  assign _0485_ = data_req_allowed_t0 & stall_ld_hz_t0;
  assign _0699_ = _0337_ | _0338_;
  assign _0700_ = _0340_ | _0341_;
  assign _0701_ = _0343_ | _0344_;
  assign _0750_ = _0438_ | _0439_;
  assign _0751_ = _0441_ | _0442_;
  assign _0752_ = _0444_ | _0445_;
  assign _0753_ = _0447_ | _0448_;
  assign _0754_ = _0450_ | _0451_;
  assign _0755_ = _0453_ | _0454_;
  assign _0756_ = _0456_ | _0457_;
  assign _0757_ = _0459_ | _0460_;
  assign _0758_ = _0462_ | _0463_;
  assign _0759_ = _0465_ | _0466_;
  assign _0760_ = _0468_ | _0469_;
  assign _0761_ = _0471_ | _0472_;
  assign _0762_ = _0474_ | _0475_;
  assign _0763_ = _0477_ | _0478_;
  assign _0764_ = _0480_ | _0481_;
  assign _0765_ = _0483_ | _0484_;
  assign _0638_ = _0699_ | _0339_;
  assign _0640_ = _0700_ | _0342_;
  assign _0642_ = _0701_ | _0345_;
  assign _0955_ = _0750_ | _0440_;
  assign multdiv_en_dec_t0 = _0751_ | _0443_;
  assign _0957_ = _0752_ | _0446_;
  assign _0959_ = _0753_ | _0449_;
  assign _0960_ = _0754_ | _0452_;
  assign _0962_ = _0755_ | _0455_;
  assign _0964_ = _0756_ | _0458_;
  assign _0966_ = _0757_ | _0461_;
  assign _0968_ = _0758_ | _0464_;
  assign stall_id_t0 = _0759_ | _0467_;
  assign _0970_ = _0760_ | _0470_;
  assign _0972_ = _0761_ | _0473_;
  assign \gen_stall_mem.instr_kill_t0  = _0762_ | _0476_;
  assign _0974_ = _0763_ | _0479_;
  assign _0976_ = _0764_ | _0482_;
  assign _0978_ = _0765_ | _0485_;
  assign _0637_ = _0981_ | _0979_;
  assign _0639_ = _0989_ | _0987_;
  assign _0641_ = _1023_ | _1021_;
  assign _0896_ = _0979_ ? _1031_ : imm_u_type;
  assign _0898_ = _0985_ ? imm_i_type : 32'd4;
  assign _0900_ = _0983_ ? imm_s_type : _0898_;
  assign imm_b = _0637_ ? _0896_ : _0900_;
  assign _0902_ = _0987_ ? imm_j_type : imm_b_type;
  assign _0904_ = _0991_ ? imm_i_type : _1031_;
  assign bt_b_operand_o = _0639_ ? _0902_ : _0904_;
  assign _0006_ = id_fsm_q ? _0056_ : _0028_;
  assign _0014_ = id_fsm_q ? 1'h0 : _0036_;
  assign _0012_ = id_fsm_q ? _0052_ : _0034_;
  assign _0018_ = id_fsm_q ? _0049_ : 1'h0;
  assign _0016_ = id_fsm_q ? _0047_ : _0038_;
  assign _0020_ = id_fsm_q ? _0054_ : _0040_;
  assign _0008_ = id_fsm_q ? 1'h0 : _0030_;
  assign _0000_ = id_fsm_q ? 1'h0 : _0022_;
  assign _0002_ = id_fsm_q ? 1'h0 : _0024_;
  assign _0010_ = id_fsm_q ? 1'h0 : _0032_;
  assign rf_wdata_id_o = rf_wdata_sel ? csr_rdata_i : result_ex_i;
  assign _0906_ = _1021_ ? imm_a : pc_id_i;
  assign _0908_ = _1025_ ? lsu_addr_last_i : multdiv_operand_a_ex_o;
  assign alu_operand_a_ex_o = _0641_ ? _0906_ : _0908_;
  assign _0184_ = | { instr_executing_spec_t0, instr_executing_t0 };
  assign _0698_ = { instr_executing, instr_executing_spec } | { instr_executing_t0, instr_executing_spec_t0 };
  assign _0183_ = & _0698_;
  assign _0092_ = _0184_ & _0183_;
  assign _0910_ = csr_op_o == 2'h1;
  assign _0912_ = csr_op_o == 2'h2;
  assign _0914_ = instr_rdata_i[31:20] == 12'h300;
  assign _0916_ = instr_rdata_i[31:20] == 12'h304;
  assign _0918_ = instr_rdata_i[31:20] == 12'h7b0;
  assign _0920_ = instr_rdata_i[31:20] == 12'h7b1;
  assign _0922_ = instr_rdata_i[31:20] == 12'h7b2;
  assign _0924_ = instr_rdata_i[31:20] == 12'h7b3;
  assign _0926_ = rf_waddr_wb_i == rf_raddr_a_o;
  assign _0928_ = rf_waddr_wb_i == rf_raddr_b_o;
  assign _0930_ = csr_op_en_o && _0934_;
  assign _0932_ = csr_op_en_o && _0942_;
  assign _0934_ = _0910_ || _0912_;
  assign _0936_ = _0914_ || _0916_;
  assign _0937_ = _0918_ || _0920_;
  assign _0939_ = _0937_ || _0922_;
  assign _0941_ = _0939_ || _0924_;
  assign _0942_ = | csr_op_o;
  assign _0944_ = ~ illegal_insn_o;
  assign _0945_ = ~ instr_valid_clear_o;
  assign _0946_ = ~ stall_id;
  assign _0947_ = ~ flush_id;
  assign _0948_ = ~ lsu_resp_valid_i;
  assign _0949_ = ~ controller_run;
  assign _0951_ = ~ ready_wb_i;
  assign _0950_ = ~ \gen_stall_mem.instr_kill ;
  assign _0952_ = ~ ebrk_insn;
  assign _0953_ = ~ ecall_insn_dec;
  assign _0954_ = illegal_insn_dec | illegal_csr_insn_i;
  assign multdiv_en_dec = mult_en_dec | div_en_dec;
  assign _0956_ = branch_set_raw | jump_set_raw;
  assign _0958_ = _0956_ | branch_jump_set_done_q;
  assign _0862_ = branch_decision_i | data_ind_timing_i;
  assign _0961_ = stall_ld_hz | stall_mem;
  assign _0963_ = _0961_ | stall_multdiv;
  assign _0965_ = _0963_ | stall_jump;
  assign _0967_ = _0965_ | stall_branch;
  assign stall_id = _0967_ | stall_alu;
  assign _0969_ = outstanding_load_wb_i | outstanding_store_wb_i;
  assign _0971_ = instr_fetch_err_i | wb_exception;
  assign \gen_stall_mem.instr_kill  = _0971_ | _0949_;
  assign _0973_ = \gen_stall_mem.outstanding_memory_access  | _0079_;
  assign _0975_ = \gen_stall_mem.rf_rd_a_hz  | \gen_stall_mem.rf_rd_b_hz ;
  assign _0977_ = \gen_stall_mem.outstanding_memory_access  | stall_ld_hz;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) branch_jump_set_done_q <= 1'h0;
    else branch_jump_set_done_q <= branch_jump_set_done_d;
  assign _0979_ = imm_b_mux_sel == 3'h5;
  assign _0981_ = imm_b_mux_sel == 3'h3;
  assign _0983_ = imm_b_mux_sel == 3'h1;
  assign _0985_ = ! imm_b_mux_sel;
  assign _0987_ = bt_b_mux_sel == 3'h4;
  assign _0989_ = bt_b_mux_sel == 3'h2;
  assign _0991_ = ! bt_b_mux_sel;
  assign bt_a_operand_o = _0993_ ? multdiv_operand_a_ex_o : pc_id_i;
  assign _0993_ = ! bt_a_mux_sel;
  assign _0056_ = _0070_ ? 1'h0 : 1'h1;
  assign _0049_ = _0070_ ? 1'h0 : jump_in_dec;
  assign _0047_ = _0070_ ? 1'h0 : branch_in_dec;
  assign _0054_ = _0070_ ? 1'h0 : multdiv_en_dec;
  assign _0052_ = multdiv_en_dec ? _0068_ : rf_we_dec;
  assign _0045_ = ex_valid_i ? rf_we_dec : 1'h0;
  assign _0051_ = ex_valid_i ? 1'h0 : 1'h1;
  assign _0044_ = lsu_req_done_i ? 1'h0 : 1'h1;
  assign _0848_ = alu_multicycle_dec ? 1'h1 : 1'h0;
  assign _0996_ = branch_in_dec ? _1033_ : _0849_;
  assign _0998_ = multdiv_en_dec ? _0051_ : _0996_;
  assign _0028_ = lsu_req_dec ? _0044_ : _0998_;
  assign _0849_ = jump_in_dec ? 1'h0 : _0848_;
  assign _0850_ = branch_in_dec ? 1'h0 : _0849_;
  assign _0851_ = multdiv_en_dec ? 1'h0 : _0850_;
  assign _0036_ = lsu_req_dec ? 1'h0 : _0851_;
  assign _1002_ = alu_multicycle_dec ? 1'h0 : rf_we_dec;
  assign _1004_ = jump_in_dec ? rf_we_dec : _1002_;
  assign _1006_ = branch_in_dec ? rf_we_dec : _1004_;
  assign _1008_ = multdiv_en_dec ? _0045_ : _1006_;
  assign _0034_ = lsu_req_dec ? rf_we_dec : _1008_;
  assign _0856_ = branch_in_dec ? data_ind_timing_i : 1'h0;
  assign _0857_ = multdiv_en_dec ? 1'h0 : _0856_;
  assign _0038_ = lsu_req_dec ? 1'h0 : _0857_;
  assign _0858_ = multdiv_en_dec ? _0051_ : 1'h0;
  assign _0040_ = lsu_req_dec ? 1'h0 : _0858_;
  assign _0859_ = jump_in_dec ? jump_set_dec : 1'h0;
  assign _0860_ = branch_in_dec ? 1'h0 : _0859_;
  assign _0861_ = multdiv_en_dec ? 1'h0 : _0860_;
  assign _0030_ = lsu_req_dec ? 1'h0 : _0861_;
  assign _0863_ = branch_in_dec ? _0862_ : 1'h0;
  assign _0864_ = multdiv_en_dec ? 1'h0 : _0863_;
  assign _0022_ = lsu_req_dec ? 1'h0 : _0864_;
  assign _0865_ = branch_in_dec ? branch_decision_i : 1'h0;
  assign _0866_ = multdiv_en_dec ? 1'h0 : _0865_;
  assign _0024_ = lsu_req_dec ? 1'h0 : _0866_;
  assign _0867_ = branch_in_dec ? 1'h1 : 1'h0;
  assign _0868_ = multdiv_en_dec ? 1'h0 : _0867_;
  assign _0032_ = lsu_req_dec ? 1'h0 : _0868_;
  assign stall_alu = instr_executing_spec ? _0014_ : 1'h0;
  assign rf_we_raw = instr_executing_spec ? _0012_ : rf_we_dec;
  assign stall_jump = instr_executing_spec ? _0018_ : 1'h0;
  assign stall_branch = instr_executing_spec ? _0016_ : 1'h0;
  assign stall_multdiv = instr_executing_spec ? _0020_ : 1'h0;
  assign jump_set_raw = instr_executing_spec ? _0008_ : 1'h0;
  assign branch_set_raw = instr_executing_spec ? _0000_ : 1'h0;
  assign branch_set_raw_spec = instr_executing_spec ? _0002_ : 1'h0;
  assign perf_branch_o = instr_executing_spec ? _0010_ : 1'h0;
  assign _0042_ = _0941_ ? 1'h1 : 1'h0;
  assign _0026_ = _0932_ ? _0042_ : 1'h0;
  assign _0004_ = _0936_ ? 1'h1 : 1'h0;
  assign csr_pipe_flush = _0930_ ? _0004_ : _0026_;
  assign _1021_ = alu_op_a_mux_sel == 2'h3;
  assign _1023_ = alu_op_a_mux_sel == 2'h2;
  assign _1025_ = alu_op_a_mux_sel == 2'h1;
  assign _1027_ = | rf_raddr_a_o;
  assign _1029_ = | rf_raddr_b_o;
  assign alu_op_a_mux_sel = lsu_addr_incr_req_i ? 2'h1 : alu_op_a_mux_sel_dec;
  assign alu_op_b_mux_sel = lsu_addr_incr_req_i ? 1'h1 : alu_op_b_mux_sel_dec;
  assign imm_b_mux_sel = lsu_addr_incr_req_i ? 3'h6 : imm_b_mux_sel_dec;
  assign imm_a = imm_a_mux_sel ? 32'd0 : zimm_rs1_type;
  assign _1031_ = instr_is_compressed_i ? 32'd2 : 32'd4;
  assign alu_operand_b_ex_o = alu_op_b_mux_sel ? imm_b : lsu_wdata_o;
  assign lsu_req_o = instr_executing ? _0064_ : 1'h0;
  assign mult_en_ex_o = instr_executing ? mult_en_dec : 1'h0;
  assign div_en_ex_o = instr_executing ? div_en_dec : 1'h0;
  assign _1033_ = data_ind_timing_i ? 1'h1 : 1'h0;
  assign multicycle_done = lsu_req_dec ? _0139_ : ex_valid_i;
  assign multdiv_operand_a_ex_o = _0081_ ? rf_wdata_fwd_wb_i : rf_rdata_a_i;
  assign lsu_wdata_o = _0083_ ? rf_wdata_fwd_wb_i : rf_rdata_b_i;
  assign _1034_ = lsu_we_o ? 2'h1 : 2'h0;
  assign instr_type_wb_o = lsu_req_dec ? _1034_ : 2'h2;
  paramodauxy_ibex_controllerWritebackStage11BranchPredictor10  controller_i (
    .branch_not_set_i(1'h0),
    .branch_not_set_i_t0(1'h0),
    .branch_set_i(branch_set),
    .branch_set_i_t0(branch_set_t0),
    .branch_set_spec_i(branch_set_spec),
    .branch_set_spec_i_t0(branch_set_spec_t0),
    .clk_i(clk_i),
    .controller_run_o(controller_run),
    .controller_run_o_t0(controller_run_t0),
    .csr_mstatus_mie_i(csr_mstatus_mie_i),
    .csr_mstatus_mie_i_t0(csr_mstatus_mie_i_t0),
    .csr_mstatus_tw_i(csr_mstatus_tw_i),
    .csr_mstatus_tw_i_t0(csr_mstatus_tw_i_t0),
    .csr_mtval_o(csr_mtval_o),
    .csr_mtval_o_t0(csr_mtval_o_t0),
    .csr_pipe_flush_i(csr_pipe_flush),
    .csr_pipe_flush_i_t0(csr_pipe_flush_t0),
    .csr_restore_dret_id_o(csr_restore_dret_id_o),
    .csr_restore_dret_id_o_t0(csr_restore_dret_id_o_t0),
    .csr_restore_mret_id_o(csr_restore_mret_id_o),
    .csr_restore_mret_id_o_t0(csr_restore_mret_id_o_t0),
    .csr_save_cause_o(csr_save_cause_o),
    .csr_save_cause_o_t0(csr_save_cause_o_t0),
    .csr_save_id_o(csr_save_id_o),
    .csr_save_id_o_t0(csr_save_id_o_t0),
    .csr_save_if_o(csr_save_if_o),
    .csr_save_if_o_t0(csr_save_if_o_t0),
    .csr_save_wb_o(csr_save_wb_o),
    .csr_save_wb_o_t0(csr_save_wb_o_t0),
    .ctrl_busy_o(ctrl_busy_o),
    .ctrl_busy_o_t0(ctrl_busy_o_t0),
    .debug_cause_o(debug_cause_o),
    .debug_cause_o_t0(debug_cause_o_t0),
    .debug_csr_save_o(debug_csr_save_o),
    .debug_csr_save_o_t0(debug_csr_save_o_t0),
    .debug_ebreakm_i(debug_ebreakm_i),
    .debug_ebreakm_i_t0(debug_ebreakm_i_t0),
    .debug_ebreaku_i(debug_ebreaku_i),
    .debug_ebreaku_i_t0(debug_ebreaku_i_t0),
    .debug_mode_o(debug_mode_o),
    .debug_mode_o_t0(debug_mode_o_t0),
    .debug_req_i(debug_req_i),
    .debug_req_i_t0(debug_req_i_t0),
    .debug_single_step_i(debug_single_step_i),
    .debug_single_step_i_t0(debug_single_step_i_t0),
    .dret_insn_i(dret_insn_dec),
    .dret_insn_i_t0(dret_insn_dec_t0),
    .ebrk_insn_i(ebrk_insn),
    .ebrk_insn_i_t0(ebrk_insn_t0),
    .ecall_insn_i(ecall_insn_dec),
    .ecall_insn_i_t0(ecall_insn_dec_t0),
    .exc_cause_o(exc_cause_o),
    .exc_cause_o_t0(exc_cause_o_t0),
    .exc_pc_mux_o(exc_pc_mux_o),
    .exc_pc_mux_o_t0(exc_pc_mux_o_t0),
    .flush_id_o(flush_id),
    .flush_id_o_t0(flush_id_t0),
    .id_in_ready_o(id_in_ready_o),
    .id_in_ready_o_t0(id_in_ready_o_t0),
    .illegal_insn_i(illegal_insn_o),
    .illegal_insn_i_t0(illegal_insn_o_t0),
    .instr_bp_taken_i(instr_bp_taken_i),
    .instr_bp_taken_i_t0(instr_bp_taken_i_t0),
    .instr_compressed_i(instr_rdata_c_i),
    .instr_compressed_i_t0(instr_rdata_c_i_t0),
    .instr_fetch_err_i(instr_fetch_err_i),
    .instr_fetch_err_i_t0(instr_fetch_err_i_t0),
    .instr_fetch_err_plus2_i(instr_fetch_err_plus2_i),
    .instr_fetch_err_plus2_i_t0(instr_fetch_err_plus2_i_t0),
    .instr_i(instr_rdata_i),
    .instr_i_t0(instr_rdata_i_t0),
    .instr_is_compressed_i(instr_is_compressed_i),
    .instr_is_compressed_i_t0(instr_is_compressed_i_t0),
    .instr_req_o(instr_req_o),
    .instr_req_o_t0(instr_req_o_t0),
    .instr_valid_clear_o(instr_valid_clear_o),
    .instr_valid_clear_o_t0(instr_valid_clear_o_t0),
    .instr_valid_i(instr_valid_i),
    .instr_valid_i_t0(instr_valid_i_t0),
    .irq_nm_i(irq_nm_i),
    .irq_nm_i_t0(irq_nm_i_t0),
    .irq_pending_i(irq_pending_i),
    .irq_pending_i_t0(irq_pending_i_t0),
    .irqs_i(irqs_i),
    .irqs_i_t0(irqs_i_t0),
    .jump_set_i(jump_set),
    .jump_set_i_t0(jump_set_t0),
    .load_err_i(lsu_load_err_i),
    .load_err_i_t0(lsu_load_err_i_t0),
    .lsu_addr_last_i(lsu_addr_last_i),
    .lsu_addr_last_i_t0(lsu_addr_last_i_t0),
    .mret_insn_i(mret_insn_dec),
    .mret_insn_i_t0(mret_insn_dec_t0),
    .nmi_mode_o(nmi_mode_o),
    .nmi_mode_o_t0(nmi_mode_o_t0),
    .nt_branch_mispredict_o(nt_branch_mispredict_o),
    .nt_branch_mispredict_o_t0(nt_branch_mispredict_o_t0),
    .pc_id_i(pc_id_i),
    .pc_id_i_t0(pc_id_i_t0),
    .pc_mux_o(pc_mux_o),
    .pc_mux_o_t0(pc_mux_o_t0),
    .pc_set_o(pc_set_o),
    .pc_set_o_t0(pc_set_o_t0),
    .pc_set_spec_o(pc_set_spec_o),
    .pc_set_spec_o_t0(pc_set_spec_o_t0),
    .perf_jump_o(perf_jump_o),
    .perf_jump_o_t0(perf_jump_o_t0),
    .perf_tbranch_o(perf_tbranch_o),
    .perf_tbranch_o_t0(perf_tbranch_o_t0),
    .priv_mode_i(priv_mode_i),
    .priv_mode_i_t0(priv_mode_i_t0),
    .ready_wb_i(ready_wb_i),
    .ready_wb_i_t0(ready_wb_i_t0),
    .rst_ni(rst_ni),
    .stall_id_i(stall_id),
    .stall_id_i_t0(stall_id_t0),
    .stall_wb_i(stall_wb),
    .stall_wb_i_t0(stall_wb_t0),
    .store_err_i(lsu_store_err_i),
    .store_err_i_t0(lsu_store_err_i_t0),
    .trigger_match_i(trigger_match_i),
    .trigger_match_i_t0(trigger_match_i_t0),
    .wb_exception_o(wb_exception),
    .wb_exception_o_t0(wb_exception_t0),
    .wfi_insn_i(wfi_insn_dec),
    .wfi_insn_i_t0(wfi_insn_dec_t0)
  );
  paramodab788080a2d62bee953947d554df7ff9d159e451auxy_ibex_decoder  decoder_i (
    .alu_multicycle_o(alu_multicycle_dec),
    .alu_multicycle_o_t0(alu_multicycle_dec_t0),
    .alu_op_a_mux_sel_o(alu_op_a_mux_sel_dec),
    .alu_op_a_mux_sel_o_t0(alu_op_a_mux_sel_dec_t0),
    .alu_op_b_mux_sel_o(alu_op_b_mux_sel_dec),
    .alu_op_b_mux_sel_o_t0(alu_op_b_mux_sel_dec_t0),
    .alu_operator_o(alu_operator_ex_o),
    .alu_operator_o_t0(alu_operator_ex_o_t0),
    .branch_in_dec_o(branch_in_dec),
    .branch_in_dec_o_t0(branch_in_dec_t0),
    .branch_taken_i(1'h1),
    .branch_taken_i_t0(1'h0),
    .bt_a_mux_sel_o(bt_a_mux_sel),
    .bt_a_mux_sel_o_t0(bt_a_mux_sel_t0),
    .bt_b_mux_sel_o(bt_b_mux_sel),
    .bt_b_mux_sel_o_t0(bt_b_mux_sel_t0),
    .clk_i(clk_i),
    .csr_access_o(csr_access_o),
    .csr_access_o_t0(csr_access_o_t0),
    .csr_op_o(csr_op_o),
    .csr_op_o_t0(csr_op_o_t0),
    .data_req_o(lsu_req_dec),
    .data_req_o_t0(lsu_req_dec_t0),
    .data_sign_extension_o(lsu_sign_ext_o),
    .data_sign_extension_o_t0(lsu_sign_ext_o_t0),
    .data_type_o(lsu_type_o),
    .data_type_o_t0(lsu_type_o_t0),
    .data_we_o(lsu_we_o),
    .data_we_o_t0(lsu_we_o_t0),
    .div_en_o(div_en_dec),
    .div_en_o_t0(div_en_dec_t0),
    .div_sel_o(div_sel_ex_o),
    .div_sel_o_t0(div_sel_ex_o_t0),
    .dret_insn_o(dret_insn_dec),
    .dret_insn_o_t0(dret_insn_dec_t0),
    .ebrk_insn_o(ebrk_insn),
    .ebrk_insn_o_t0(ebrk_insn_t0),
    .ecall_insn_o(ecall_insn_dec),
    .ecall_insn_o_t0(ecall_insn_dec_t0),
    .icache_inval_o(icache_inval_o),
    .icache_inval_o_t0(icache_inval_o_t0),
    .illegal_c_insn_i(illegal_c_insn_i),
    .illegal_c_insn_i_t0(illegal_c_insn_i_t0),
    .illegal_insn_o(illegal_insn_dec),
    .illegal_insn_o_t0(illegal_insn_dec_t0),
    .imm_a_mux_sel_o(imm_a_mux_sel),
    .imm_a_mux_sel_o_t0(imm_a_mux_sel_t0),
    .imm_b_mux_sel_o(imm_b_mux_sel_dec),
    .imm_b_mux_sel_o_t0(imm_b_mux_sel_dec_t0),
    .imm_b_type_o(imm_b_type),
    .imm_b_type_o_t0(imm_b_type_t0),
    .imm_i_type_o(imm_i_type),
    .imm_i_type_o_t0(imm_i_type_t0),
    .imm_j_type_o(imm_j_type),
    .imm_j_type_o_t0(imm_j_type_t0),
    .imm_s_type_o(imm_s_type),
    .imm_s_type_o_t0(imm_s_type_t0),
    .imm_u_type_o(imm_u_type),
    .imm_u_type_o_t0(imm_u_type_t0),
    .instr_first_cycle_i(instr_first_cycle_id_o),
    .instr_first_cycle_i_t0(instr_first_cycle_id_o_t0),
    .instr_rdata_alu_i(instr_rdata_alu_i),
    .instr_rdata_alu_i_t0(instr_rdata_alu_i_t0),
    .instr_rdata_i(instr_rdata_i),
    .instr_rdata_i_t0(instr_rdata_i_t0),
    .jump_in_dec_o(jump_in_dec),
    .jump_in_dec_o_t0(jump_in_dec_t0),
    .jump_set_o(jump_set_dec),
    .jump_set_o_t0(jump_set_dec_t0),
    .mret_insn_o(mret_insn_dec),
    .mret_insn_o_t0(mret_insn_dec_t0),
    .mult_en_o(mult_en_dec),
    .mult_en_o_t0(mult_en_dec_t0),
    .mult_sel_o(mult_sel_ex_o),
    .mult_sel_o_t0(mult_sel_ex_o_t0),
    .multdiv_operator_o(multdiv_operator_ex_o),
    .multdiv_operator_o_t0(multdiv_operator_ex_o_t0),
    .multdiv_signed_mode_o(multdiv_signed_mode_ex_o),
    .multdiv_signed_mode_o_t0(multdiv_signed_mode_ex_o_t0),
    .rf_raddr_a_o(rf_raddr_a_o),
    .rf_raddr_a_o_t0(rf_raddr_a_o_t0),
    .rf_raddr_b_o(rf_raddr_b_o),
    .rf_raddr_b_o_t0(rf_raddr_b_o_t0),
    .rf_ren_a_o(rf_ren_a_dec),
    .rf_ren_a_o_t0(rf_ren_a_dec_t0),
    .rf_ren_b_o(rf_ren_b_dec),
    .rf_ren_b_o_t0(rf_ren_b_dec_t0),
    .rf_waddr_o(rf_waddr_id_o),
    .rf_waddr_o_t0(rf_waddr_id_o_t0),
    .rf_wdata_sel_o(rf_wdata_sel),
    .rf_wdata_sel_o_t0(rf_wdata_sel_t0),
    .rf_we_o(rf_we_dec),
    .rf_we_o_t0(rf_we_dec_t0),
    .rst_ni(rst_ni),
    .wfi_insn_o(wfi_insn_dec),
    .wfi_insn_o_t0(wfi_insn_dec_t0),
    .zimm_rs1_type_o(zimm_rs1_type),
    .zimm_rs1_type_o_t0(zimm_rs1_type_t0)
  );
  assign multdiv_operand_b_ex_o = lsu_wdata_o;
  assign multdiv_operand_b_ex_o_t0 = lsu_wdata_o_t0;
  assign multdiv_ready_id_o = ready_wb_i;
  assign multdiv_ready_id_o_t0 = ready_wb_i_t0;
endmodule

module paramodeccb28a0d9c7c379466a9299a8885e9ec9033585auxy_ibex_csr (clk_i, rst_ni, wr_data_i, wr_en_i, rd_data_o, rd_error_o, rd_data_o_t0, rd_error_o_t0, wr_data_i_t0, wr_en_i_t0);
  wire _00_;
  wire _01_;
  wire _02_;
  wire _03_;
  wire _04_;
  wire _05_;
  wire _06_;
  wire _07_;
  wire _08_;
  input clk_i;
  wire clk_i;
  output rd_data_o;
  reg rd_data_o;
  output rd_data_o_t0;
  reg rd_data_o_t0;
  output rd_error_o;
  wire rd_error_o;
  output rd_error_o_t0;
  wire rd_error_o_t0;
  input rst_ni;
  wire rst_ni;
  input wr_data_i;
  wire wr_data_i;
  input wr_data_i_t0;
  wire wr_data_i_t0;
  input wr_en_i;
  wire wr_en_i;
  input wr_en_i_t0;
  wire wr_en_i_t0;
  assign _00_ = ~ wr_en_i;
  assign _08_ = wr_data_i ^ rd_data_o;
  assign _04_ = wr_data_i_t0 | rd_data_o_t0;
  assign _05_ = _08_ | _04_;
  assign _01_ = wr_en_i & wr_data_i_t0;
  assign _02_ = _00_ & rd_data_o_t0;
  assign _03_ = _05_ & wr_en_i_t0;
  assign _06_ = _01_ | _02_;
  assign _07_ = _06_ | _03_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) rd_data_o_t0 <= 1'h0;
    else rd_data_o_t0 <= _07_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) rd_data_o <= 1'h0;
    else if (wr_en_i) rd_data_o <= wr_data_i;
  assign rd_error_o = 1'h0;
  assign rd_error_o_t0 = 1'h0;
endmodule

module paramodauxy_ibex_aluRV32Bs3200000000000000000000000000000000 (operator_i, operand_a_i, operand_b_i, instr_first_cycle_i, multdiv_operand_a_i, multdiv_operand_b_i, multdiv_sel_i, imd_val_q_i, imd_val_d_o, imd_val_we_o, adder_result_o, adder_result_ext_o, result_o, comparison_result_o, is_equal_result_o, instr_first_cycle_i_t0, adder_result_ext_o_t0, adder_result_o_t0, comparison_result_o_t0, imd_val_d_o_t0, imd_val_q_i_t0
, imd_val_we_o_t0, is_equal_result_o_t0, multdiv_operand_a_i_t0, multdiv_operand_b_i_t0, multdiv_sel_i_t0, operand_a_i_t0, operand_b_i_t0, operator_i_t0, result_o_t0);
  wire _0000_;
  wire _0001_;
  wire [33:0] _0002_;
  wire [33:0] _0003_;
  wire _0004_;
  wire _0005_;
  wire _0006_;
  wire _0007_;
  wire [31:0] _0008_;
  wire [31:0] _0009_;
  wire [31:0] _0010_;
  wire [31:0] _0011_;
  wire _0012_;
  wire _0013_;
  wire [31:0] _0014_;
  wire _0015_;
  wire _0016_;
  wire _0017_;
  wire _0018_;
  wire _0019_;
  wire [31:0] _0020_;
  wire [31:0] _0021_;
  wire _0022_;
  wire _0023_;
  wire _0024_;
  wire _0025_;
  wire [7:0] _0026_;
  wire [5:0] _0027_;
  wire [4:0] _0028_;
  wire [1:0] _0029_;
  wire [5:0] _0030_;
  wire [31:0] _0031_;
  wire [31:0] _0032_;
  wire [5:0] _0033_;
  wire [3:0] _0034_;
  wire _0035_;
  wire [4:0] _0036_;
  wire [32:0] _0037_;
  wire [32:0] _0038_;
  wire [5:0] _0039_;
  wire [31:0] _0040_;
  wire [4:0] _0041_;
  wire [31:0] _0042_;
  wire _0043_;
  wire _0044_;
  wire _0045_;
  wire _0046_;
  wire _0047_;
  wire _0048_;
  wire _0049_;
  wire _0050_;
  wire _0051_;
  wire _0052_;
  wire _0053_;
  wire _0054_;
  wire _0055_;
  wire _0056_;
  wire _0057_;
  wire _0058_;
  wire _0059_;
  wire _0060_;
  wire _0061_;
  wire _0062_;
  wire [33:0] _0063_;
  wire [33:0] _0064_;
  wire _0065_;
  wire _0066_;
  wire _0067_;
  wire [31:0] _0068_;
  wire [31:0] _0069_;
  wire [31:0] _0070_;
  wire _0071_;
  wire _0072_;
  wire _0073_;
  wire _0074_;
  wire _0075_;
  wire _0076_;
  wire [31:0] _0077_;
  wire [31:0] _0078_;
  wire [31:0] _0079_;
  wire [31:0] _0080_;
  wire [31:0] _0081_;
  wire [31:0] _0082_;
  wire [31:0] _0083_;
  wire [31:0] _0084_;
  wire [31:0] _0085_;
  wire [31:0] _0086_;
  wire [31:0] _0087_;
  wire [31:0] _0088_;
  wire _0089_;
  wire _0090_;
  wire _0091_;
  wire _0092_;
  wire _0093_;
  wire _0094_;
  wire _0095_;
  wire _0096_;
  wire _0097_;
  wire [31:0] _0098_;
  wire _0099_;
  wire _0100_;
  wire _0101_;
  wire _0102_;
  wire _0103_;
  wire _0104_;
  wire _0105_;
  wire _0106_;
  wire _0107_;
  wire _0108_;
  wire _0109_;
  wire _0110_;
  wire _0111_;
  wire _0112_;
  wire _0113_;
  wire _0114_;
  wire _0115_;
  wire _0116_;
  wire _0117_;
  wire _0118_;
  wire _0119_;
  wire _0120_;
  wire _0121_;
  wire _0122_;
  wire _0123_;
  wire _0124_;
  wire _0125_;
  wire _0126_;
  wire [31:0] _0127_;
  wire [31:0] _0128_;
  wire _0129_;
  wire _0130_;
  wire _0131_;
  wire _0132_;
  wire _0133_;
  wire _0134_;
  wire [7:0] _0135_;
  wire [5:0] _0136_;
  wire [5:0] _0137_;
  wire [4:0] _0138_;
  wire [5:0] _0139_;
  wire [5:0] _0140_;
  wire [5:0] _0141_;
  wire [5:0] _0142_;
  wire [1:0] _0143_;
  wire [5:0] _0144_;
  wire [5:0] _0145_;
  wire [5:0] _0146_;
  wire [5:0] _0147_;
  wire [5:0] _0148_;
  wire [5:0] _0149_;
  wire [5:0] _0150_;
  wire [5:0] _0151_;
  wire [31:0] _0152_;
  wire [31:0] _0153_;
  wire [31:0] _0154_;
  wire [31:0] _0155_;
  wire [31:0] _0156_;
  wire [31:0] _0157_;
  wire [5:0] _0158_;
  wire [5:0] _0159_;
  wire [5:0] _0160_;
  wire [5:0] _0161_;
  wire [5:0] _0162_;
  wire [5:0] _0163_;
  wire [5:0] _0164_;
  wire [5:0] _0165_;
  wire [3:0] _0166_;
  wire [5:0] _0167_;
  wire [5:0] _0168_;
  wire [5:0] _0169_;
  wire [5:0] _0170_;
  wire [5:0] _0171_;
  wire _0172_;
  wire _0173_;
  wire _0174_;
  wire [4:0] _0175_;
  wire [32:0] _0176_;
  wire [32:0] _0177_;
  wire [32:0] _0178_;
  wire [32:0] _0179_;
  wire [32:0] _0180_;
  wire [32:0] _0181_;
  wire [5:0] _0182_;
  wire [5:0] _0183_;
  wire [5:0] _0184_;
  wire [5:0] _0185_;
  wire [5:0] _0186_;
  wire [5:0] _0187_;
  wire [5:0] _0188_;
  wire [5:0] _0189_;
  wire [5:0] _0190_;
  wire [5:0] _0191_;
  wire [5:0] _0192_;
  wire [5:0] _0193_;
  wire [5:0] _0194_;
  wire [5:0] _0195_;
  wire [5:0] _0196_;
  wire [5:0] _0197_;
  wire [5:0] _0198_;
  wire [5:0] _0199_;
  wire [5:0] _0200_;
  wire [5:0] _0201_;
  wire [5:0] _0202_;
  wire [5:0] _0203_;
  wire [5:0] _0204_;
  wire [5:0] _0205_;
  wire [5:0] _0206_;
  wire [5:0] _0207_;
  wire [5:0] _0208_;
  wire [5:0] _0209_;
  wire [5:0] _0210_;
  wire [5:0] _0211_;
  wire [5:0] _0212_;
  wire [5:0] _0213_;
  wire [527:0] _0214_;
  wire [32:0] _0215_;
  wire [31:0] _0216_;
  wire [4:0] _0217_;
  wire [4:0] _0218_;
  wire [4:0] _0219_;
  wire [31:0] _0220_;
  wire [31:0] _0221_;
  wire [31:0] _0222_;
  wire [31:0] _0223_;
  wire [31:0] _0224_;
  wire [31:0] _0225_;
  wire [32:0] _0226_;
  wire [32:0] _0227_;
  wire [32:0] _0228_;
  wire _0229_;
  wire _0230_;
  wire _0231_;
  wire _0232_;
  wire [33:0] _0233_;
  wire [33:0] _0234_;
  wire [33:0] _0235_;
  wire _0236_;
  wire [31:0] _0237_;
  wire _0238_;
  wire _0239_;
  wire [31:0] _0240_;
  wire [31:0] _0241_;
  wire [31:0] _0242_;
  wire [31:0] _0243_;
  wire [31:0] _0244_;
  wire [31:0] _0245_;
  wire [31:0] _0246_;
  wire [31:0] _0247_;
  wire [31:0] _0248_;
  wire [31:0] _0249_;
  wire [31:0] _0250_;
  wire [31:0] _0251_;
  wire _0252_;
  wire _0253_;
  wire _0254_;
  wire _0255_;
  wire _0256_;
  wire _0257_;
  wire _0258_;
  wire _0259_;
  wire _0260_;
  wire _0261_;
  wire _0262_;
  wire _0263_;
  wire _0264_;
  wire _0265_;
  wire _0266_;
  wire _0267_;
  wire _0268_;
  wire _0269_;
  wire _0270_;
  wire _0271_;
  wire _0272_;
  wire _0273_;
  wire _0274_;
  wire [31:0] _0275_;
  wire _0276_;
  wire _0277_;
  wire [31:0] _0278_;
  wire [31:0] _0279_;
  wire [31:0] _0280_;
  wire [31:0] _0281_;
  wire [31:0] _0282_;
  wire [31:0] _0283_;
  wire _0284_;
  wire _0285_;
  wire _0286_;
  wire [32:0] _0287_;
  wire [32:0] _0288_;
  wire [32:0] _0289_;
  wire [32:0] _0290_;
  wire [32:0] _0291_;
  wire [32:0] _0292_;
  wire [527:0] _0293_;
  wire [527:0] _0294_;
  wire [32:0] _0295_;
  wire [31:0] _0296_;
  wire [31:0] _0297_;
  wire [4:0] _0298_;
  wire [4:0] _0299_;
  wire [4:0] _0300_;
  wire [31:0] _0301_;
  wire [31:0] _0302_;
  wire [31:0] _0303_;
  wire [31:0] _0304_;
  wire [32:0] _0305_;
  wire [33:0] _0306_;
  wire [31:0] _0307_;
  wire [31:0] _0308_;
  wire [31:0] _0309_;
  wire _0310_;
  wire _0311_;
  wire _0312_;
  wire _0313_;
  wire _0314_;
  wire _0315_;
  wire _0316_;
  wire _0317_;
  wire _0318_;
  wire _0319_;
  wire _0320_;
  wire _0321_;
  wire _0322_;
  wire _0323_;
  wire [31:0] _0324_;
  wire [31:0] _0325_;
  wire _0326_;
  wire [32:0] _0327_;
  wire [32:0] _0328_;
  wire [527:0] _0329_;
  wire [32:0] _0330_;
  wire [4:0] _0331_;
  wire [31:0] _0332_;
  wire [31:0] _0333_;
  wire [32:0] _0334_;
  wire _0335_;
  wire _0336_;
  wire _0337_;
  wire _0338_;
  wire _0339_;
  wire _0340_;
  wire _0341_;
  wire _0342_;
  wire _0343_;
  wire _0344_;
  wire _0345_;
  wire _0346_;
  wire _0347_;
  wire _0348_;
  wire _0349_;
  wire _0350_;
  wire _0351_;
  wire _0352_;
  wire _0353_;
  wire _0354_;
  wire _0355_;
  wire _0356_;
  wire _0357_;
  wire _0358_;
  wire _0359_;
  wire _0360_;
  wire _0361_;
  wire _0362_;
  wire _0363_;
  wire _0364_;
  wire _0365_;
  wire _0366_;
  wire _0367_;
  wire _0368_;
  wire _0369_;
  wire _0370_;
  wire _0371_;
  wire _0372_;
  wire _0373_;
  wire _0374_;
  wire _0375_;
  wire _0376_;
  wire _0377_;
  wire _0378_;
  wire _0379_;
  wire _0380_;
  wire _0381_;
  wire _0382_;
  wire _0383_;
  wire _0384_;
  wire _0385_;
  wire _0386_;
  wire _0387_;
  wire _0388_;
  wire _0389_;
  wire _0390_;
  wire _0391_;
  wire _0392_;
  wire _0393_;
  wire _0394_;
  wire _0395_;
  wire _0396_;
  wire _0397_;
  wire _0398_;
  wire _0399_;
  wire _0400_;
  wire _0401_;
  wire _0402_;
  wire _0403_;
  wire _0404_;
  wire _0405_;
  wire _0406_;
  wire _0407_;
  wire _0408_;
  wire _0409_;
  wire _0410_;
  wire _0411_;
  wire _0412_;
  wire _0413_;
  wire _0414_;
  wire _0415_;
  wire _0416_;
  wire _0417_;
  wire _0418_;
  wire _0419_;
  wire _0420_;
  wire _0421_;
  wire _0422_;
  wire [33:0] _0423_;
  wire [33:0] _0424_;
  wire [31:0] _0425_;
  wire [31:0] _0426_;
  wire [31:0] _0427_;
  wire [31:0] _0428_;
  wire [31:0] _0429_;
  wire [31:0] _0430_;
  wire [31:0] _0431_;
  wire [31:0] _0432_;
  wire _0433_;
  wire _0434_;
  wire _0435_;
  wire _0436_;
  wire [32:0] _0437_;
  wire [32:0] _0438_;
  wire _0439_;
  wire _0440_;
  wire _0441_;
  wire _0442_;
  wire _0443_;
  wire _0444_;
  wire _0445_;
  wire _0446_;
  wire _0447_;
  wire _0448_;
  wire _0449_;
  wire _0450_;
  wire _0451_;
  wire _0452_;
  wire _0453_;
  wire _0454_;
  wire _0455_;
  wire _0456_;
  wire _0457_;
  wire _0458_;
  wire _0459_;
  wire _0460_;
  wire _0461_;
  wire _0462_;
  wire _0463_;
  wire _0464_;
  wire _0465_;
  wire _0466_;
  wire _0467_;
  wire _0468_;
  wire _0469_;
  wire _0470_;
  wire [7:0] _0471_;
  wire [7:0] _0472_;
  wire _0473_;
  wire _0474_;
  wire [4:0] _0475_;
  wire [4:0] _0476_;
  wire _0477_;
  wire _0478_;
  wire [1:0] _0479_;
  wire [1:0] _0480_;
  wire _0481_;
  wire _0482_;
  wire [5:0] _0483_;
  wire [5:0] _0484_;
  wire _0485_;
  wire _0486_;
  wire [31:0] _0487_;
  wire [31:0] _0488_;
  wire [5:0] _0489_;
  wire [5:0] _0490_;
  wire _0491_;
  wire _0492_;
  wire [3:0] _0493_;
  wire [3:0] _0494_;
  wire _0495_;
  wire _0496_;
  wire _0497_;
  wire [32:0] _0498_;
  wire [32:0] _0499_;
  wire [31:0] _0500_;
  wire [31:0] _0501_;
  wire _0502_;
  wire _0503_;
  wire _0504_;
  wire _0505_;
  wire [32:0] adder_in_a;
  wire [32:0] adder_in_a_t0;
  wire [32:0] adder_in_b;
  wire [32:0] adder_in_b_t0;
  wire adder_op_b_negate;
  wire adder_op_b_negate_t0;
  output [33:0] adder_result_ext_o;
  wire [33:0] adder_result_ext_o;
  output [33:0] adder_result_ext_o_t0;
  wire [33:0] adder_result_ext_o_t0;
  output [31:0] adder_result_o;
  wire [31:0] adder_result_o;
  output [31:0] adder_result_o_t0;
  wire [31:0] adder_result_o_t0;
  wire bwlogic_and;
  wire [31:0] bwlogic_and_result;
  wire [31:0] bwlogic_and_result_t0;
  wire bwlogic_and_t0;
  wire bwlogic_or;
  wire [31:0] bwlogic_or_result;
  wire [31:0] bwlogic_or_result_t0;
  wire bwlogic_or_t0;
  wire [31:0] bwlogic_result;
  wire [31:0] bwlogic_result_t0;
  wire [31:0] bwlogic_xor_result;
  wire [31:0] bwlogic_xor_result_t0;
  wire cmp_signed;
  wire cmp_signed_t0;
  output comparison_result_o;
  wire comparison_result_o;
  output comparison_result_o_t0;
  wire comparison_result_o_t0;
  output [63:0] imd_val_d_o;
  wire [63:0] imd_val_d_o;
  output [63:0] imd_val_d_o_t0;
  wire [63:0] imd_val_d_o_t0;
  input [63:0] imd_val_q_i;
  wire [63:0] imd_val_q_i;
  input [63:0] imd_val_q_i_t0;
  wire [63:0] imd_val_q_i_t0;
  output [1:0] imd_val_we_o;
  wire [1:0] imd_val_we_o;
  output [1:0] imd_val_we_o_t0;
  wire [1:0] imd_val_we_o_t0;
  input instr_first_cycle_i;
  wire instr_first_cycle_i;
  input instr_first_cycle_i_t0;
  wire instr_first_cycle_i_t0;
  output is_equal_result_o;
  wire is_equal_result_o;
  output is_equal_result_o_t0;
  wire is_equal_result_o_t0;
  wire is_greater_equal;
  wire is_greater_equal_t0;
  input [32:0] multdiv_operand_a_i;
  wire [32:0] multdiv_operand_a_i;
  input [32:0] multdiv_operand_a_i_t0;
  wire [32:0] multdiv_operand_a_i_t0;
  input [32:0] multdiv_operand_b_i;
  wire [32:0] multdiv_operand_b_i;
  input [32:0] multdiv_operand_b_i_t0;
  wire [32:0] multdiv_operand_b_i_t0;
  input multdiv_sel_i;
  wire multdiv_sel_i;
  input multdiv_sel_i_t0;
  wire multdiv_sel_i_t0;
  input [31:0] operand_a_i;
  wire [31:0] operand_a_i;
  input [31:0] operand_a_i_t0;
  wire [31:0] operand_a_i_t0;
  input [31:0] operand_b_i;
  wire [31:0] operand_b_i;
  input [31:0] operand_b_i_t0;
  wire [31:0] operand_b_i_t0;
  wire [32:0] operand_b_neg;
  input [5:0] operator_i;
  wire [5:0] operator_i;
  input [5:0] operator_i_t0;
  wire [5:0] operator_i_t0;
  output [31:0] result_o;
  wire [31:0] result_o;
  output [31:0] result_o_t0;
  wire [31:0] result_o_t0;
  wire [5:0] shift_amt;
  wire [5:0] shift_amt_compl;
  wire [5:0] shift_amt_compl_t0;
  wire [5:0] shift_amt_t0;
  wire shift_arith;
  wire shift_arith_t0;
  wire shift_left;
  wire shift_left_t0;
  wire [31:0] shift_operand;
  wire [31:0] shift_operand_t0;
  wire [31:0] shift_result;
  wire [32:0] shift_result_ext;
  wire [32:0] shift_result_ext_t0;
  wire [31:0] shift_result_t0;
  assign adder_result_ext_o = { 1'h0, adder_in_a } + { 1'h0, adder_in_b };
  assign _0000_ = shift_arith & shift_operand[31];
  assign bwlogic_and_result = operand_a_i & operand_b_i;
  assign _0002_ = ~ { 1'h0, adder_in_a_t0 };
  assign _0003_ = ~ { 1'h0, adder_in_b_t0 };
  assign _0063_ = { 1'h0, adder_in_a } & _0002_;
  assign _0064_ = { 1'h0, adder_in_b } & _0003_;
  assign _0423_ = _0063_ + _0064_;
  assign _0233_ = { 1'h0, adder_in_a } | { 1'h0, adder_in_a_t0 };
  assign _0234_ = { 1'h0, adder_in_b } | { 1'h0, adder_in_b_t0 };
  assign _0424_ = _0233_ + _0234_;
  assign _0306_ = _0423_ ^ _0424_;
  assign _0235_ = _0306_ | { 1'h0, adder_in_a_t0 };
  assign adder_result_ext_o_t0 = _0235_ | { 1'h0, adder_in_b_t0 };
  assign _0065_ = shift_arith_t0 & shift_operand[31];
  assign _0068_ = operand_a_i_t0 & operand_b_i;
  assign _0066_ = shift_operand_t0[31] & shift_arith;
  assign _0069_ = operand_b_i_t0 & operand_a_i;
  assign _0067_ = shift_arith_t0 & shift_operand_t0[31];
  assign _0236_ = _0065_ | _0066_;
  assign _0237_ = _0068_ | _0069_;
  assign _0001_ = _0236_ | _0067_;
  assign bwlogic_and_result_t0 = _0237_ | _0070_;
  assign _0047_ = | operator_i_t0;
  assign _0027_ = ~ operator_i_t0;
  assign _0136_ = operator_i & _0027_;
  assign _0137_ = 6'h17 & _0027_;
  assign _0139_ = 6'h09 & _0027_;
  assign _0140_ = 6'h08 & _0027_;
  assign _0141_ = 6'h0c & _0027_;
  assign _0142_ = 6'h0b & _0027_;
  assign _0144_ = 6'h01 & _0027_;
  assign _0146_ = 6'h02 & _0027_;
  assign _0147_ = 6'h05 & _0027_;
  assign _0148_ = 6'h03 & _0027_;
  assign _0149_ = 6'h06 & _0027_;
  assign _0150_ = 6'h04 & _0027_;
  assign _0151_ = 6'h07 & _0027_;
  assign _0158_ = 6'h0a & _0027_;
  assign _0160_ = 6'h13 & _0027_;
  assign _0161_ = 6'h14 & _0027_;
  assign _0162_ = 6'h19 & _0027_;
  assign _0163_ = 6'h1a & _0027_;
  assign _0164_ = 6'h25 & _0027_;
  assign _0165_ = 6'h26 & _0027_;
  assign _0167_ = 6'h15 & _0027_;
  assign _0168_ = 6'h16 & _0027_;
  assign _0169_ = 6'h1b & _0027_;
  assign _0170_ = 6'h1c & _0027_;
  assign _0171_ = 6'h18 & _0027_;
  assign _0335_ = _0136_ == _0137_;
  assign _0336_ = _0136_ == _0139_;
  assign _0337_ = _0136_ == _0140_;
  assign _0338_ = _0136_ == _0141_;
  assign _0339_ = _0136_ == _0142_;
  assign _0340_ = _0136_ == _0144_;
  assign _0341_ = _0136_ == _0146_;
  assign _0342_ = _0136_ == _0147_;
  assign _0343_ = _0136_ == _0148_;
  assign _0344_ = _0136_ == _0149_;
  assign _0345_ = _0136_ == _0150_;
  assign _0346_ = _0136_ == _0151_;
  assign _0347_ = _0136_ == _0158_;
  assign _0348_ = _0136_ == _0160_;
  assign _0349_ = _0136_ == _0161_;
  assign _0350_ = _0136_ == _0162_;
  assign _0351_ = _0136_ == _0163_;
  assign _0352_ = _0136_ == _0164_;
  assign _0353_ = _0136_ == _0165_;
  assign _0354_ = _0136_ == _0167_;
  assign _0355_ = _0136_ == _0168_;
  assign _0356_ = _0136_ == _0169_;
  assign _0357_ = _0136_ == _0170_;
  assign _0358_ = _0136_ == _0171_;
  assign _0472_[0] = _0335_ & _0047_;
  assign _0476_[1] = _0336_ & _0047_;
  assign shift_arith_t0 = _0337_ & _0047_;
  assign _0476_[3] = _0338_ & _0047_;
  assign _0476_[4] = _0339_ & _0047_;
  assign _0480_[1] = _0340_ & _0047_;
  assign _0484_[0] = _0341_ & _0047_;
  assign _0484_[1] = _0342_ & _0047_;
  assign _0440_ = _0343_ & _0047_;
  assign _0442_ = _0344_ & _0047_;
  assign _0444_ = _0345_ & _0047_;
  assign _0446_ = _0346_ & _0047_;
  assign shift_left_t0 = _0347_ & _0047_;
  assign _0472_[4] = _0348_ & _0047_;
  assign _0472_[5] = _0349_ & _0047_;
  assign _0490_[2] = _0350_ & _0047_;
  assign _0490_[3] = _0351_ & _0047_;
  assign _0472_[6] = _0352_ & _0047_;
  assign _0472_[7] = _0353_ & _0047_;
  assign _0472_[2] = _0354_ & _0047_;
  assign _0472_[3] = _0355_ & _0047_;
  assign _0494_[2] = _0356_ & _0047_;
  assign _0494_[3] = _0357_ & _0047_;
  assign _0472_[1] = _0358_ & _0047_;
  assign _0045_ = | adder_result_ext_o_t0[32:1];
  assign _0046_ = | _0472_;
  assign _0048_ = | { shift_left_t0, _0476_[4:3], _0476_[1], shift_arith_t0 };
  assign _0049_ = | _0480_;
  assign _0050_ = | { _0484_[1:0], _0446_, _0444_, _0442_, _0440_ };
  assign _0051_ = | { _0490_[3:2], _0472_[7:4] };
  assign _0052_ = | { _0494_[3:2], _0472_[3:2] };
  assign _0053_ = | { _0494_[2], _0490_[2], _0472_[6], _0472_[4], _0472_[2] };
  assign _0014_ = ~ adder_result_ext_o_t0[32:1];
  assign _0026_ = ~ _0472_;
  assign _0028_ = ~ { _0476_[4:3], _0476_[1], shift_left_t0, shift_arith_t0 };
  assign _0029_ = ~ _0480_;
  assign _0030_ = ~ { _0484_[1:0], _0446_, _0444_, _0442_, _0440_ };
  assign _0033_ = ~ { _0490_[3:2], _0472_[7:4] };
  assign _0034_ = ~ { _0494_[3:2], _0472_[3:2] };
  assign _0036_ = ~ { _0494_[2], _0490_[2], _0472_[6], _0472_[4], _0472_[2] };
  assign _0098_ = adder_result_ext_o[32:1] & _0014_;
  assign _0135_ = _0471_ & _0026_;
  assign _0138_ = { _0475_[4:3], _0475_[1:0], shift_arith } & _0028_;
  assign _0143_ = _0479_ & _0029_;
  assign _0145_ = { _0483_[1:0], _0445_, _0443_, _0441_, _0439_ } & _0030_;
  assign _0159_ = { _0489_[3:2], _0471_[7:4] } & _0033_;
  assign _0166_ = { _0493_[3:2], _0471_[3:2] } & _0034_;
  assign _0175_ = { _0493_[2], _0489_[2], _0471_[6], _0471_[4], _0471_[2] } & _0036_;
  assign _0054_ = ! _0098_;
  assign _0055_ = ! _0135_;
  assign _0056_ = ! _0138_;
  assign _0057_ = ! _0143_;
  assign _0058_ = ! _0136_;
  assign _0059_ = ! _0145_;
  assign _0060_ = ! _0159_;
  assign _0061_ = ! _0166_;
  assign _0062_ = ! _0175_;
  assign is_equal_result_o_t0 = _0054_ & _0045_;
  assign _0474_ = _0055_ & _0046_;
  assign _0478_ = _0056_ & _0048_;
  assign _0482_ = _0057_ & _0049_;
  assign _0480_[0] = _0058_ & _0047_;
  assign _0486_ = _0059_ & _0050_;
  assign _0492_ = _0060_ & _0051_;
  assign _0496_ = _0061_ & _0052_;
  assign cmp_signed_t0 = _0062_ & _0053_;
  assign _0008_ = ~ { _0473_, _0473_, _0473_, _0473_, _0473_, _0473_, _0473_, _0473_, _0473_, _0473_, _0473_, _0473_, _0473_, _0473_, _0473_, _0473_, _0473_, _0473_, _0473_, _0473_, _0473_, _0473_, _0473_, _0473_, _0473_, _0473_, _0473_, _0473_, _0473_, _0473_, _0473_, _0473_ };
  assign _0009_ = ~ { _0485_, _0485_, _0485_, _0485_, _0485_, _0485_, _0485_, _0485_, _0485_, _0485_, _0485_, _0485_, _0485_, _0485_, _0485_, _0485_, _0485_, _0485_, _0485_, _0485_, _0485_, _0485_, _0485_, _0485_, _0485_, _0485_, _0485_, _0485_, _0485_, _0485_, _0485_, _0485_ };
  assign _0010_ = ~ { _0481_, _0481_, _0481_, _0481_, _0481_, _0481_, _0481_, _0481_, _0481_, _0481_, _0481_, _0481_, _0481_, _0481_, _0481_, _0481_, _0481_, _0481_, _0481_, _0481_, _0481_, _0481_, _0481_, _0481_, _0481_, _0481_, _0481_, _0481_, _0481_, _0481_, _0481_, _0481_ };
  assign _0011_ = ~ { _0229_, _0229_, _0229_, _0229_, _0229_, _0229_, _0229_, _0229_, _0229_, _0229_, _0229_, _0229_, _0229_, _0229_, _0229_, _0229_, _0229_, _0229_, _0229_, _0229_, _0229_, _0229_, _0229_, _0229_, _0229_, _0229_, _0229_, _0229_, _0229_, _0229_, _0229_, _0229_ };
  assign _0007_ = ~ _0491_;
  assign _0012_ = ~ _0471_[1];
  assign _0013_ = ~ _0231_;
  assign _0015_ = ~ operator_i[5];
  assign _0016_ = ~ operator_i[4];
  assign _0017_ = ~ operator_i[3];
  assign _0018_ = ~ operator_i[2];
  assign _0019_ = ~ operator_i[1];
  assign _0031_ = ~ { bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and };
  assign _0032_ = ~ { bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or };
  assign _0035_ = ~ _0502_;
  assign _0037_ = ~ { adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate };
  assign _0038_ = ~ { multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i };
  assign _0041_ = ~ { instr_first_cycle_i, instr_first_cycle_i, instr_first_cycle_i, instr_first_cycle_i, instr_first_cycle_i };
  assign _0042_ = ~ { shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left };
  assign _0240_ = { _0474_, _0474_, _0474_, _0474_, _0474_, _0474_, _0474_, _0474_, _0474_, _0474_, _0474_, _0474_, _0474_, _0474_, _0474_, _0474_, _0474_, _0474_, _0474_, _0474_, _0474_, _0474_, _0474_, _0474_, _0474_, _0474_, _0474_, _0474_, _0474_, _0474_, _0474_, _0474_ } | _0008_;
  assign _0243_ = { _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_ } | _0009_;
  assign _0246_ = { _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_ } | _0010_;
  assign _0249_ = { _0230_, _0230_, _0230_, _0230_, _0230_, _0230_, _0230_, _0230_, _0230_, _0230_, _0230_, _0230_, _0230_, _0230_, _0230_, _0230_, _0230_, _0230_, _0230_, _0230_, _0230_, _0230_, _0230_, _0230_, _0230_, _0230_, _0230_, _0230_, _0230_, _0230_, _0230_, _0230_ } | _0011_;
  assign _0252_ = _0492_ | _0007_;
  assign _0255_ = _0472_[1] | _0012_;
  assign _0258_ = _0232_ | _0013_;
  assign _0261_ = operator_i_t0[5] | _0015_;
  assign _0264_ = operator_i_t0[4] | _0016_;
  assign _0267_ = operator_i_t0[3] | _0017_;
  assign _0270_ = operator_i_t0[2] | _0018_;
  assign _0272_ = operator_i_t0[1] | _0019_;
  assign _0278_ = { bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0 } | _0031_;
  assign _0281_ = { bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0 } | _0032_;
  assign _0284_ = _0503_ | _0035_;
  assign _0287_ = { adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0 } | _0037_;
  assign _0290_ = { multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0 } | _0038_;
  assign _0298_ = { instr_first_cycle_i_t0, instr_first_cycle_i_t0, instr_first_cycle_i_t0, instr_first_cycle_i_t0, instr_first_cycle_i_t0 } | _0041_;
  assign _0301_ = { shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0 } | _0042_;
  assign _0241_ = { _0474_, _0474_, _0474_, _0474_, _0474_, _0474_, _0474_, _0474_, _0474_, _0474_, _0474_, _0474_, _0474_, _0474_, _0474_, _0474_, _0474_, _0474_, _0474_, _0474_, _0474_, _0474_, _0474_, _0474_, _0474_, _0474_, _0474_, _0474_, _0474_, _0474_, _0474_, _0474_ } | { _0473_, _0473_, _0473_, _0473_, _0473_, _0473_, _0473_, _0473_, _0473_, _0473_, _0473_, _0473_, _0473_, _0473_, _0473_, _0473_, _0473_, _0473_, _0473_, _0473_, _0473_, _0473_, _0473_, _0473_, _0473_, _0473_, _0473_, _0473_, _0473_, _0473_, _0473_, _0473_ };
  assign _0244_ = { _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_ } | { _0485_, _0485_, _0485_, _0485_, _0485_, _0485_, _0485_, _0485_, _0485_, _0485_, _0485_, _0485_, _0485_, _0485_, _0485_, _0485_, _0485_, _0485_, _0485_, _0485_, _0485_, _0485_, _0485_, _0485_, _0485_, _0485_, _0485_, _0485_, _0485_, _0485_, _0485_, _0485_ };
  assign _0247_ = { _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_ } | { _0481_, _0481_, _0481_, _0481_, _0481_, _0481_, _0481_, _0481_, _0481_, _0481_, _0481_, _0481_, _0481_, _0481_, _0481_, _0481_, _0481_, _0481_, _0481_, _0481_, _0481_, _0481_, _0481_, _0481_, _0481_, _0481_, _0481_, _0481_, _0481_, _0481_, _0481_, _0481_ };
  assign _0250_ = { _0230_, _0230_, _0230_, _0230_, _0230_, _0230_, _0230_, _0230_, _0230_, _0230_, _0230_, _0230_, _0230_, _0230_, _0230_, _0230_, _0230_, _0230_, _0230_, _0230_, _0230_, _0230_, _0230_, _0230_, _0230_, _0230_, _0230_, _0230_, _0230_, _0230_, _0230_, _0230_ } | { _0229_, _0229_, _0229_, _0229_, _0229_, _0229_, _0229_, _0229_, _0229_, _0229_, _0229_, _0229_, _0229_, _0229_, _0229_, _0229_, _0229_, _0229_, _0229_, _0229_, _0229_, _0229_, _0229_, _0229_, _0229_, _0229_, _0229_, _0229_, _0229_, _0229_, _0229_, _0229_ };
  assign _0253_ = _0492_ | _0491_;
  assign _0256_ = _0472_[1] | _0471_[1];
  assign _0259_ = _0232_ | _0231_;
  assign _0262_ = operator_i_t0[5] | operator_i[5];
  assign _0265_ = operator_i_t0[4] | operator_i[4];
  assign _0268_ = operator_i_t0[3] | operator_i[3];
  assign _0271_ = operator_i_t0[2] | operator_i[2];
  assign _0273_ = operator_i_t0[1] | operator_i[1];
  assign _0279_ = { bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0 } | { bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and };
  assign _0282_ = { bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0 } | { bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or };
  assign _0285_ = _0503_ | _0502_;
  assign _0288_ = { adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0 } | { adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate };
  assign _0291_ = { multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0 } | { multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i };
  assign _0299_ = { instr_first_cycle_i_t0, instr_first_cycle_i_t0, instr_first_cycle_i_t0, instr_first_cycle_i_t0, instr_first_cycle_i_t0 } | { instr_first_cycle_i, instr_first_cycle_i, instr_first_cycle_i, instr_first_cycle_i, instr_first_cycle_i };
  assign _0302_ = { shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0 } | { shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left };
  assign _0077_ = shift_result_t0 & _0240_;
  assign _0080_ = 32'd0 & _0243_;
  assign _0083_ = _0430_ & _0246_;
  assign _0086_ = _0432_ & _0249_;
  assign _0089_ = is_greater_equal_t0 & _0252_;
  assign _0092_ = is_equal_result_o_t0 & _0255_;
  assign _0095_ = _0436_ & _0258_;
  assign _0099_ = _0449_ & _0261_;
  assign _0102_ = _0453_ & _0264_;
  assign _0105_ = _0456_ & _0264_;
  assign _0107_ = _0457_ & _0267_;
  assign _0109_ = _0459_ & _0267_;
  assign _0112_ = _0462_ & _0267_;
  assign _0114_ = _0463_ & _0270_;
  assign _0116_ = _0465_ & _0270_;
  assign _0122_ = operator_i_t0[0] & _0272_;
  assign _0152_ = bwlogic_xor_result_t0 & _0278_;
  assign _0155_ = _0488_ & _0281_;
  assign _0172_ = adder_result_ext_o_t0[32] & _0284_;
  assign _0176_ = { operand_b_i_t0, 1'h0 } & _0287_;
  assign _0179_ = _0499_ & _0290_;
  assign _0217_ = shift_amt_compl_t0[4:0] & _0298_;
  assign _0220_ = operand_a_i_t0 & _0301_;
  assign _0223_ = shift_result_ext_t0[31:0] & _0301_;
  assign _0226_ = { operand_a_i_t0, 1'h0 } & _0290_;
  assign _0078_ = { 31'h00000000, comparison_result_o_t0 } & _0241_;
  assign _0081_ = bwlogic_result_t0 & _0244_;
  assign _0084_ = adder_result_ext_o_t0[32:1] & _0247_;
  assign _0087_ = _0428_ & _0250_;
  assign _0090_ = is_greater_equal_t0 & _0253_;
  assign _0093_ = is_equal_result_o_t0 & _0256_;
  assign _0096_ = _0434_ & _0259_;
  assign _0100_ = _0451_ & _0262_;
  assign _0103_ = _0455_ & _0265_;
  assign _0110_ = _0461_ & _0268_;
  assign _0118_ = _0467_ & _0271_;
  assign _0120_ = _0468_ & _0271_;
  assign _0124_ = operator_i_t0[0] & _0273_;
  assign _0153_ = bwlogic_and_result_t0 & _0279_;
  assign _0156_ = bwlogic_or_result_t0 & _0282_;
  assign _0173_ = _0505_ & _0285_;
  assign _0177_ = { operand_b_i_t0, 1'h0 } & _0288_;
  assign _0180_ = multdiv_operand_b_i_t0 & _0291_;
  assign _0218_ = operand_b_i_t0[4:0] & _0299_;
  assign _0221_ = { operand_a_i_t0[0], operand_a_i_t0[1], operand_a_i_t0[2], operand_a_i_t0[3], operand_a_i_t0[4], operand_a_i_t0[5], operand_a_i_t0[6], operand_a_i_t0[7], operand_a_i_t0[8], operand_a_i_t0[9], operand_a_i_t0[10], operand_a_i_t0[11], operand_a_i_t0[12], operand_a_i_t0[13], operand_a_i_t0[14], operand_a_i_t0[15], operand_a_i_t0[16], operand_a_i_t0[17], operand_a_i_t0[18], operand_a_i_t0[19], operand_a_i_t0[20], operand_a_i_t0[21], operand_a_i_t0[22], operand_a_i_t0[23], operand_a_i_t0[24], operand_a_i_t0[25], operand_a_i_t0[26], operand_a_i_t0[27], operand_a_i_t0[28], operand_a_i_t0[29], operand_a_i_t0[30], operand_a_i_t0[31] } & _0302_;
  assign _0224_ = { shift_result_ext_t0[0], shift_result_ext_t0[1], shift_result_ext_t0[2], shift_result_ext_t0[3], shift_result_ext_t0[4], shift_result_ext_t0[5], shift_result_ext_t0[6], shift_result_ext_t0[7], shift_result_ext_t0[8], shift_result_ext_t0[9], shift_result_ext_t0[10], shift_result_ext_t0[11], shift_result_ext_t0[12], shift_result_ext_t0[13], shift_result_ext_t0[14], shift_result_ext_t0[15], shift_result_ext_t0[16], shift_result_ext_t0[17], shift_result_ext_t0[18], shift_result_ext_t0[19], shift_result_ext_t0[20], shift_result_ext_t0[21], shift_result_ext_t0[22], shift_result_ext_t0[23], shift_result_ext_t0[24], shift_result_ext_t0[25], shift_result_ext_t0[26], shift_result_ext_t0[27], shift_result_ext_t0[28], shift_result_ext_t0[29], shift_result_ext_t0[30], shift_result_ext_t0[31] } & _0302_;
  assign _0227_ = multdiv_operand_a_i_t0 & _0291_;
  assign _0242_ = _0077_ | _0078_;
  assign _0245_ = _0080_ | _0081_;
  assign _0248_ = _0083_ | _0084_;
  assign _0251_ = _0086_ | _0087_;
  assign _0254_ = _0089_ | _0090_;
  assign _0257_ = _0092_ | _0093_;
  assign _0260_ = _0095_ | _0096_;
  assign _0263_ = _0099_ | _0100_;
  assign _0266_ = _0102_ | _0103_;
  assign _0269_ = _0109_ | _0110_;
  assign _0274_ = _0122_ | _0124_;
  assign _0280_ = _0152_ | _0153_;
  assign _0283_ = _0155_ | _0156_;
  assign _0286_ = _0172_ | _0173_;
  assign _0289_ = _0176_ | _0177_;
  assign _0292_ = _0179_ | _0180_;
  assign _0300_ = _0217_ | _0218_;
  assign _0303_ = _0220_ | _0221_;
  assign _0304_ = _0223_ | _0224_;
  assign _0305_ = _0226_ | _0227_;
  assign _0307_ = shift_result ^ { 31'h00000000, comparison_result_o };
  assign _0308_ = _0429_ ^ adder_result_ext_o[32:1];
  assign _0309_ = _0431_ ^ _0427_;
  assign _0310_ = is_greater_equal ^ _0470_;
  assign _0311_ = is_equal_result_o ^ _0469_;
  assign _0312_ = _0435_ ^ _0433_;
  assign _0313_ = _0448_ ^ _0450_;
  assign _0314_ = _0452_ ^ _0454_;
  assign _0317_ = _0458_ ^ _0460_;
  assign _0323_ = _0321_ ^ _0322_;
  assign _0324_ = bwlogic_xor_result ^ bwlogic_and_result;
  assign _0325_ = _0487_ ^ bwlogic_or_result;
  assign _0326_ = _0447_ ^ _0504_;
  assign _0327_ = { operand_b_i, 1'h0 } ^ operand_b_neg;
  assign _0328_ = _0498_ ^ multdiv_operand_b_i;
  assign _0331_ = shift_amt_compl[4:0] ^ operand_b_i[4:0];
  assign _0332_ = operand_a_i ^ { operand_a_i[0], operand_a_i[1], operand_a_i[2], operand_a_i[3], operand_a_i[4], operand_a_i[5], operand_a_i[6], operand_a_i[7], operand_a_i[8], operand_a_i[9], operand_a_i[10], operand_a_i[11], operand_a_i[12], operand_a_i[13], operand_a_i[14], operand_a_i[15], operand_a_i[16], operand_a_i[17], operand_a_i[18], operand_a_i[19], operand_a_i[20], operand_a_i[21], operand_a_i[22], operand_a_i[23], operand_a_i[24], operand_a_i[25], operand_a_i[26], operand_a_i[27], operand_a_i[28], operand_a_i[29], operand_a_i[30], operand_a_i[31] };
  assign _0333_ = shift_result_ext[31:0] ^ { shift_result_ext[0], shift_result_ext[1], shift_result_ext[2], shift_result_ext[3], shift_result_ext[4], shift_result_ext[5], shift_result_ext[6], shift_result_ext[7], shift_result_ext[8], shift_result_ext[9], shift_result_ext[10], shift_result_ext[11], shift_result_ext[12], shift_result_ext[13], shift_result_ext[14], shift_result_ext[15], shift_result_ext[16], shift_result_ext[17], shift_result_ext[18], shift_result_ext[19], shift_result_ext[20], shift_result_ext[21], shift_result_ext[22], shift_result_ext[23], shift_result_ext[24], shift_result_ext[25], shift_result_ext[26], shift_result_ext[27], shift_result_ext[28], shift_result_ext[29], shift_result_ext[30], shift_result_ext[31] };
  assign _0334_ = { operand_a_i, 1'h1 } ^ multdiv_operand_a_i;
  assign _0079_ = { _0474_, _0474_, _0474_, _0474_, _0474_, _0474_, _0474_, _0474_, _0474_, _0474_, _0474_, _0474_, _0474_, _0474_, _0474_, _0474_, _0474_, _0474_, _0474_, _0474_, _0474_, _0474_, _0474_, _0474_, _0474_, _0474_, _0474_, _0474_, _0474_, _0474_, _0474_, _0474_ } & _0307_;
  assign _0082_ = { _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_ } & bwlogic_result;
  assign _0085_ = { _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_ } & _0308_;
  assign _0088_ = { _0230_, _0230_, _0230_, _0230_, _0230_, _0230_, _0230_, _0230_, _0230_, _0230_, _0230_, _0230_, _0230_, _0230_, _0230_, _0230_, _0230_, _0230_, _0230_, _0230_, _0230_, _0230_, _0230_, _0230_, _0230_, _0230_, _0230_, _0230_, _0230_, _0230_, _0230_, _0230_ } & _0309_;
  assign _0091_ = _0492_ & _0310_;
  assign _0094_ = _0472_[1] & _0311_;
  assign _0097_ = _0232_ & _0312_;
  assign _0101_ = operator_i_t0[5] & _0313_;
  assign _0104_ = operator_i_t0[4] & _0314_;
  assign _0106_ = operator_i_t0[4] & _0315_;
  assign _0108_ = operator_i_t0[3] & _0316_;
  assign _0111_ = operator_i_t0[3] & _0317_;
  assign _0113_ = operator_i_t0[3] & _0318_;
  assign _0115_ = operator_i_t0[2] & _0319_;
  assign _0117_ = operator_i_t0[2] & _0043_;
  assign _0119_ = operator_i_t0[2] & _0044_;
  assign _0121_ = operator_i_t0[2] & _0320_;
  assign _0123_ = operator_i_t0[1] & _0321_;
  assign _0125_ = operator_i_t0[1] & _0322_;
  assign _0126_ = operator_i_t0[1] & _0323_;
  assign _0154_ = { bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0 } & _0324_;
  assign _0157_ = { bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0 } & _0325_;
  assign _0174_ = _0503_ & _0326_;
  assign _0178_ = { adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0 } & _0327_;
  assign _0181_ = { multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0 } & _0328_;
  assign _0219_ = { instr_first_cycle_i_t0, instr_first_cycle_i_t0, instr_first_cycle_i_t0, instr_first_cycle_i_t0, instr_first_cycle_i_t0 } & _0331_;
  assign _0222_ = { shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0 } & _0332_;
  assign _0225_ = { shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0 } & _0333_;
  assign _0228_ = { multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0 } & _0334_;
  assign _0428_ = _0079_ | _0242_;
  assign _0430_ = _0082_ | _0245_;
  assign _0432_ = _0085_ | _0248_;
  assign result_o_t0 = _0088_ | _0251_;
  assign _0434_ = _0091_ | _0254_;
  assign _0436_ = _0094_ | _0257_;
  assign comparison_result_o_t0 = _0097_ | _0260_;
  assign adder_op_b_negate_t0 = _0101_ | _0263_;
  assign _0449_ = _0104_ | _0266_;
  assign _0451_ = _0106_ | _0105_;
  assign _0453_ = _0108_ | _0107_;
  assign _0455_ = _0111_ | _0269_;
  assign _0456_ = _0113_ | _0112_;
  assign _0457_ = _0115_ | _0114_;
  assign _0459_ = _0117_ | _0116_;
  assign _0461_ = _0119_ | _0118_;
  assign _0462_ = _0121_ | _0120_;
  assign _0463_ = _0123_ | _0122_;
  assign _0465_ = _0123_ | _0124_;
  assign _0467_ = _0125_ | _0122_;
  assign _0468_ = _0126_ | _0274_;
  assign _0488_ = _0154_ | _0280_;
  assign bwlogic_result_t0 = _0157_ | _0283_;
  assign is_greater_equal_t0 = _0174_ | _0286_;
  assign _0499_ = _0178_ | _0289_;
  assign adder_in_b_t0 = _0181_ | _0292_;
  assign shift_amt_t0[4:0] = _0219_ | _0300_;
  assign shift_operand_t0 = _0222_ | _0303_;
  assign shift_result_t0 = _0225_ | _0304_;
  assign adder_in_a_t0 = _0228_ | _0305_;
  assign _0043_ = ~ _0464_;
  assign _0044_ = ~ _0466_;
  assign _0004_ = ~ _0477_;
  assign _0006_ = ~ _0495_;
  assign _0020_ = ~ operand_a_i;
  assign _0022_ = ~ _0439_;
  assign _0024_ = ~ _0443_;
  assign _0005_ = ~ _0473_;
  assign _0021_ = ~ operand_b_i;
  assign _0023_ = ~ _0441_;
  assign _0025_ = ~ _0445_;
  assign _0071_ = _0478_ & _0005_;
  assign _0074_ = _0496_ & _0007_;
  assign _0127_ = operand_a_i_t0 & _0021_;
  assign _0129_ = _0440_ & _0023_;
  assign _0132_ = _0444_ & _0025_;
  assign _0072_ = _0474_ & _0004_;
  assign _0075_ = _0492_ & _0006_;
  assign _0128_ = operand_b_i_t0 & _0020_;
  assign _0130_ = _0442_ & _0022_;
  assign _0133_ = _0446_ & _0024_;
  assign _0073_ = _0478_ & _0474_;
  assign _0076_ = _0496_ & _0492_;
  assign _0070_ = operand_a_i_t0 & operand_b_i_t0;
  assign _0131_ = _0440_ & _0442_;
  assign _0134_ = _0444_ & _0446_;
  assign _0238_ = _0071_ | _0072_;
  assign _0239_ = _0074_ | _0075_;
  assign _0275_ = _0127_ | _0128_;
  assign _0276_ = _0129_ | _0130_;
  assign _0277_ = _0132_ | _0133_;
  assign _0230_ = _0238_ | _0073_;
  assign _0232_ = _0239_ | _0076_;
  assign bwlogic_or_result_t0 = _0275_ | _0070_;
  assign bwlogic_or_t0 = _0276_ | _0131_;
  assign bwlogic_and_t0 = _0277_ | _0134_;
  assign _0229_ = _0477_ | _0473_;
  assign _0231_ = _0495_ | _0491_;
  assign _0427_ = _0473_ ? { 31'h00000000, comparison_result_o } : shift_result;
  assign _0429_ = _0485_ ? bwlogic_result : 32'd0;
  assign _0431_ = _0481_ ? adder_result_ext_o[32:1] : _0429_;
  assign result_o = _0229_ ? _0427_ : _0431_;
  assign _0433_ = _0491_ ? _0470_ : is_greater_equal;
  assign _0435_ = _0471_[1] ? _0469_ : is_equal_result_o;
  assign comparison_result_o = _0231_ ? _0433_ : _0435_;
  assign _0183_ = { 1'h0, shift_amt_t0[4:0] } & 6'h01;
  assign _0184_ = { 1'h0, shift_amt_t0[4:0] } & 6'h02;
  assign _0185_ = { 1'h0, shift_amt_t0[4:0] } & 6'h03;
  assign _0186_ = { 1'h0, shift_amt_t0[4:0] } & 6'h04;
  assign _0187_ = { 1'h0, shift_amt_t0[4:0] } & 6'h05;
  assign _0188_ = { 1'h0, shift_amt_t0[4:0] } & 6'h06;
  assign _0189_ = { 1'h0, shift_amt_t0[4:0] } & 6'h07;
  assign _0190_ = { 1'h0, shift_amt_t0[4:0] } & 6'h08;
  assign _0191_ = { 1'h0, shift_amt_t0[4:0] } & 6'h09;
  assign _0192_ = { 1'h0, shift_amt_t0[4:0] } & 6'h0a;
  assign _0193_ = { 1'h0, shift_amt_t0[4:0] } & 6'h0b;
  assign _0194_ = { 1'h0, shift_amt_t0[4:0] } & 6'h0c;
  assign _0195_ = { 1'h0, shift_amt_t0[4:0] } & 6'h0d;
  assign _0196_ = { 1'h0, shift_amt_t0[4:0] } & 6'h0e;
  assign _0197_ = { 1'h0, shift_amt_t0[4:0] } & 6'h0f;
  assign _0198_ = { 1'h0, shift_amt_t0[4:0] } & 6'h10;
  assign _0199_ = { 1'h0, shift_amt_t0[4:0] } & 6'h11;
  assign _0200_ = { 1'h0, shift_amt_t0[4:0] } & 6'h12;
  assign _0201_ = { 1'h0, shift_amt_t0[4:0] } & 6'h13;
  assign _0202_ = { 1'h0, shift_amt_t0[4:0] } & 6'h14;
  assign _0203_ = { 1'h0, shift_amt_t0[4:0] } & 6'h15;
  assign _0204_ = { 1'h0, shift_amt_t0[4:0] } & 6'h16;
  assign _0205_ = { 1'h0, shift_amt_t0[4:0] } & 6'h17;
  assign _0206_ = { 1'h0, shift_amt_t0[4:0] } & 6'h18;
  assign _0207_ = { 1'h0, shift_amt_t0[4:0] } & 6'h19;
  assign _0208_ = { 1'h0, shift_amt_t0[4:0] } & 6'h1a;
  assign _0209_ = { 1'h0, shift_amt_t0[4:0] } & 6'h1b;
  assign _0210_ = { 1'h0, shift_amt_t0[4:0] } & 6'h1c;
  assign _0211_ = { 1'h0, shift_amt_t0[4:0] } & 6'h1d;
  assign _0212_ = { 1'h0, shift_amt_t0[4:0] } & 6'h1e;
  assign _0213_ = { 1'h0, shift_amt_t0[4:0] } & 6'h1f;
  assign _0359_ = _0183_ == 6'h01;
  assign _0360_ = _0184_ == 6'h02;
  assign _0361_ = _0185_ == 6'h03;
  assign _0362_ = _0186_ == 6'h04;
  assign _0363_ = _0187_ == 6'h05;
  assign _0364_ = _0188_ == 6'h06;
  assign _0365_ = _0189_ == 6'h07;
  assign _0366_ = _0190_ == 6'h08;
  assign _0367_ = _0191_ == 6'h09;
  assign _0368_ = _0192_ == 6'h0a;
  assign _0369_ = _0193_ == 6'h0b;
  assign _0370_ = _0194_ == 6'h0c;
  assign _0371_ = _0195_ == 6'h0d;
  assign _0372_ = _0196_ == 6'h0e;
  assign _0373_ = _0197_ == 6'h0f;
  assign _0374_ = _0198_ == 6'h10;
  assign _0375_ = _0199_ == 6'h11;
  assign _0376_ = _0200_ == 6'h12;
  assign _0377_ = _0201_ == 6'h13;
  assign _0378_ = _0202_ == 6'h14;
  assign _0379_ = _0203_ == 6'h15;
  assign _0380_ = _0204_ == 6'h16;
  assign _0381_ = _0205_ == 6'h17;
  assign _0382_ = _0206_ == 6'h18;
  assign _0383_ = _0207_ == 6'h19;
  assign _0384_ = _0208_ == 6'h1a;
  assign _0385_ = _0209_ == 6'h1b;
  assign _0386_ = _0210_ == 6'h1c;
  assign _0387_ = _0211_ == 6'h1d;
  assign _0388_ = _0212_ == 6'h1e;
  assign _0389_ = _0213_ == 6'h1f;
  assign _0329_ = { _0437_[31:30], _0437_[30:29], _0437_[29], _0437_[29:28], _0437_[28], _0437_[28], _0437_[28:27], _0437_[27], _0437_[27], _0437_[27], _0437_[27:26], _0437_[26], _0437_[26], _0437_[26], _0437_[26], _0437_[26:25], _0437_[25], _0437_[25], _0437_[25], _0437_[25], _0437_[25], _0437_[25:24], _0437_[24], _0437_[24], _0437_[24], _0437_[24], _0437_[24], _0437_[24], _0437_[24:23], _0437_[23], _0437_[23], _0437_[23], _0437_[23], _0437_[23], _0437_[23], _0437_[23], _0437_[23:22], _0437_[22], _0437_[22], _0437_[22], _0437_[22], _0437_[22], _0437_[22], _0437_[22], _0437_[22], _0437_[22:21], _0437_[21], _0437_[21], _0437_[21], _0437_[21], _0437_[21], _0437_[21], _0437_[21], _0437_[21], _0437_[21], _0437_[21:20], _0437_[20], _0437_[20], _0437_[20], _0437_[20], _0437_[20], _0437_[20], _0437_[20], _0437_[20], _0437_[20], _0437_[20], _0437_[20:19], _0437_[19], _0437_[19], _0437_[19], _0437_[19], _0437_[19], _0437_[19], _0437_[19], _0437_[19], _0437_[19], _0437_[19], _0437_[19], _0437_[19:18], _0437_[18], _0437_[18], _0437_[18], _0437_[18], _0437_[18], _0437_[18], _0437_[18], _0437_[18], _0437_[18], _0437_[18], _0437_[18], _0437_[18], _0437_[18:17], _0437_[17], _0437_[17], _0437_[17], _0437_[17], _0437_[17], _0437_[17], _0437_[17], _0437_[17], _0437_[17], _0437_[17], _0437_[17], _0437_[17], _0437_[17], _0437_[17:16], _0437_[16], _0437_[16], _0437_[16], _0437_[16], _0437_[16], _0437_[16], _0437_[16], _0437_[16], _0437_[16], _0437_[16], _0437_[16], _0437_[16], _0437_[16], _0437_[16], _0437_[16:15], _0437_[15], _0437_[15], _0437_[15], _0437_[15], _0437_[15], _0437_[15], _0437_[15], _0437_[15], _0437_[15], _0437_[15], _0437_[15], _0437_[15], _0437_[15], _0437_[15], _0437_[15], _0437_[15:14], _0437_[14], _0437_[14], _0437_[14], _0437_[14], _0437_[14], _0437_[14], _0437_[14], _0437_[14], _0437_[14], _0437_[14], _0437_[14], _0437_[14], _0437_[14], _0437_[14], _0437_[14], _0437_[14], _0437_[14:13], _0437_[13], _0437_[13], _0437_[13], _0437_[13], _0437_[13], _0437_[13], _0437_[13], _0437_[13], _0437_[13], _0437_[13], _0437_[13], _0437_[13], _0437_[13], _0437_[13], _0437_[13], _0437_[13], _0437_[13], _0437_[13:12], _0437_[12], _0437_[12], _0437_[12], _0437_[12], _0437_[12], _0437_[12], _0437_[12], _0437_[12], _0437_[12], _0437_[12], _0437_[12], _0437_[12], _0437_[12], _0437_[12], _0437_[12], _0437_[12], _0437_[12], _0437_[12], _0437_[12:11], _0437_[11], _0437_[11], _0437_[11], _0437_[11], _0437_[11], _0437_[11], _0437_[11], _0437_[11], _0437_[11], _0437_[11], _0437_[11], _0437_[11], _0437_[11], _0437_[11], _0437_[11], _0437_[11], _0437_[11], _0437_[11], _0437_[11], _0437_[11:10], _0437_[10], _0437_[10], _0437_[10], _0437_[10], _0437_[10], _0437_[10], _0437_[10], _0437_[10], _0437_[10], _0437_[10], _0437_[10], _0437_[10], _0437_[10], _0437_[10], _0437_[10], _0437_[10], _0437_[10], _0437_[10], _0437_[10], _0437_[10], _0437_[10:9], _0437_[9], _0437_[9], _0437_[9], _0437_[9], _0437_[9], _0437_[9], _0437_[9], _0437_[9], _0437_[9], _0437_[9], _0437_[9], _0437_[9], _0437_[9], _0437_[9], _0437_[9], _0437_[9], _0437_[9], _0437_[9], _0437_[9], _0437_[9], _0437_[9], _0437_[9:8], _0437_[8], _0437_[8], _0437_[8], _0437_[8], _0437_[8], _0437_[8], _0437_[8], _0437_[8], _0437_[8], _0437_[8], _0437_[8], _0437_[8], _0437_[8], _0437_[8], _0437_[8], _0437_[8], _0437_[8], _0437_[8], _0437_[8], _0437_[8], _0437_[8], _0437_[8], _0437_[8:7], _0437_[7], _0437_[7], _0437_[7], _0437_[7], _0437_[7], _0437_[7], _0437_[7], _0437_[7], _0437_[7], _0437_[7], _0437_[7], _0437_[7], _0437_[7], _0437_[7], _0437_[7], _0437_[7], _0437_[7], _0437_[7], _0437_[7], _0437_[7], _0437_[7], _0437_[7], _0437_[7], _0437_[7:6], _0437_[6], _0437_[6], _0437_[6], _0437_[6], _0437_[6], _0437_[6], _0437_[6], _0437_[6], _0437_[6], _0437_[6], _0437_[6], _0437_[6], _0437_[6], _0437_[6], _0437_[6], _0437_[6], _0437_[6], _0437_[6], _0437_[6], _0437_[6], _0437_[6], _0437_[6], _0437_[6], _0437_[6], _0437_[6:5], _0437_[5], _0437_[5], _0437_[5], _0437_[5], _0437_[5], _0437_[5], _0437_[5], _0437_[5], _0437_[5], _0437_[5], _0437_[5], _0437_[5], _0437_[5], _0437_[5], _0437_[5], _0437_[5], _0437_[5], _0437_[5], _0437_[5], _0437_[5], _0437_[5], _0437_[5], _0437_[5], _0437_[5], _0437_[5], _0437_[5:4], _0437_[4], _0437_[4], _0437_[4], _0437_[4], _0437_[4], _0437_[4], _0437_[4], _0437_[4], _0437_[4], _0437_[4], _0437_[4], _0437_[4], _0437_[4], _0437_[4], _0437_[4], _0437_[4], _0437_[4], _0437_[4], _0437_[4], _0437_[4], _0437_[4], _0437_[4], _0437_[4], _0437_[4], _0437_[4], _0437_[4], _0437_[4:3], _0437_[3], _0437_[3], _0437_[3], _0437_[3], _0437_[3], _0437_[3], _0437_[3], _0437_[3], _0437_[3], _0437_[3], _0437_[3], _0437_[3], _0437_[3], _0437_[3], _0437_[3], _0437_[3], _0437_[3], _0437_[3], _0437_[3], _0437_[3], _0437_[3], _0437_[3], _0437_[3], _0437_[3], _0437_[3], _0437_[3], _0437_[3], _0437_[3:2], _0437_[2], _0437_[2], _0437_[2], _0437_[2], _0437_[2], _0437_[2], _0437_[2], _0437_[2], _0437_[2], _0437_[2], _0437_[2], _0437_[2], _0437_[2], _0437_[2], _0437_[2], _0437_[2], _0437_[2], _0437_[2], _0437_[2], _0437_[2], _0437_[2], _0437_[2], _0437_[2], _0437_[2], _0437_[2], _0437_[2], _0437_[2], _0437_[2], _0437_[2:1], _0437_[1], _0437_[1], _0437_[1], _0437_[1], _0437_[1], _0437_[1], _0437_[1], _0437_[1], _0437_[1], _0437_[1], _0437_[1], _0437_[1], _0437_[1], _0437_[1], _0437_[1], _0437_[1], _0437_[1], _0437_[1], _0437_[1], _0437_[1], _0437_[1], _0437_[1], _0437_[1], _0437_[1], _0437_[1], _0437_[1], _0437_[1], _0437_[1], _0437_[1], _0437_[1:0], _0437_[0], _0437_[0], _0437_[0], _0437_[0], _0437_[0], _0437_[0], _0437_[0], _0437_[0], _0437_[0], _0437_[0], _0437_[0], _0437_[0], _0437_[0], _0437_[0], _0437_[0], _0437_[0], _0437_[0], _0437_[0], _0437_[0], _0437_[0], _0437_[0], _0437_[0], _0437_[0], _0437_[0], _0437_[0], _0437_[0], _0437_[0], _0437_[0], _0437_[0], _0437_[0], _0437_[0] } ^ { _0437_[32], _0437_[32:31], _0437_[32:30], _0437_[32:29], _0437_[32:28], _0437_[32:27], _0437_[32:26], _0437_[32:25], _0437_[32:24], _0437_[32:23], _0437_[32:22], _0437_[32:21], _0437_[32:20], _0437_[32:19], _0437_[32:18], _0437_[32:17], _0437_[32:16], _0437_[32:15], _0437_[32:14], _0437_[32:13], _0437_[32:12], _0437_[32:11], _0437_[32:10], _0437_[32:9], _0437_[32:8], _0437_[32:7], _0437_[32:6], _0437_[32:5], _0437_[32:4], _0437_[32:3], _0437_[32:2], _0437_[32:1] };
  assign _0293_ = { _0438_[31:30], _0438_[30:29], _0438_[29], _0438_[29:28], _0438_[28], _0438_[28], _0438_[28:27], _0438_[27], _0438_[27], _0438_[27], _0438_[27:26], _0438_[26], _0438_[26], _0438_[26], _0438_[26], _0438_[26:25], _0438_[25], _0438_[25], _0438_[25], _0438_[25], _0438_[25], _0438_[25:24], _0438_[24], _0438_[24], _0438_[24], _0438_[24], _0438_[24], _0438_[24], _0438_[24:23], _0438_[23], _0438_[23], _0438_[23], _0438_[23], _0438_[23], _0438_[23], _0438_[23], _0438_[23:22], _0438_[22], _0438_[22], _0438_[22], _0438_[22], _0438_[22], _0438_[22], _0438_[22], _0438_[22], _0438_[22:21], _0438_[21], _0438_[21], _0438_[21], _0438_[21], _0438_[21], _0438_[21], _0438_[21], _0438_[21], _0438_[21], _0438_[21:20], _0438_[20], _0438_[20], _0438_[20], _0438_[20], _0438_[20], _0438_[20], _0438_[20], _0438_[20], _0438_[20], _0438_[20], _0438_[20:19], _0438_[19], _0438_[19], _0438_[19], _0438_[19], _0438_[19], _0438_[19], _0438_[19], _0438_[19], _0438_[19], _0438_[19], _0438_[19], _0438_[19:18], _0438_[18], _0438_[18], _0438_[18], _0438_[18], _0438_[18], _0438_[18], _0438_[18], _0438_[18], _0438_[18], _0438_[18], _0438_[18], _0438_[18], _0438_[18:17], _0438_[17], _0438_[17], _0438_[17], _0438_[17], _0438_[17], _0438_[17], _0438_[17], _0438_[17], _0438_[17], _0438_[17], _0438_[17], _0438_[17], _0438_[17], _0438_[17:16], _0438_[16], _0438_[16], _0438_[16], _0438_[16], _0438_[16], _0438_[16], _0438_[16], _0438_[16], _0438_[16], _0438_[16], _0438_[16], _0438_[16], _0438_[16], _0438_[16], _0438_[16:15], _0438_[15], _0438_[15], _0438_[15], _0438_[15], _0438_[15], _0438_[15], _0438_[15], _0438_[15], _0438_[15], _0438_[15], _0438_[15], _0438_[15], _0438_[15], _0438_[15], _0438_[15], _0438_[15:14], _0438_[14], _0438_[14], _0438_[14], _0438_[14], _0438_[14], _0438_[14], _0438_[14], _0438_[14], _0438_[14], _0438_[14], _0438_[14], _0438_[14], _0438_[14], _0438_[14], _0438_[14], _0438_[14], _0438_[14:13], _0438_[13], _0438_[13], _0438_[13], _0438_[13], _0438_[13], _0438_[13], _0438_[13], _0438_[13], _0438_[13], _0438_[13], _0438_[13], _0438_[13], _0438_[13], _0438_[13], _0438_[13], _0438_[13], _0438_[13], _0438_[13:12], _0438_[12], _0438_[12], _0438_[12], _0438_[12], _0438_[12], _0438_[12], _0438_[12], _0438_[12], _0438_[12], _0438_[12], _0438_[12], _0438_[12], _0438_[12], _0438_[12], _0438_[12], _0438_[12], _0438_[12], _0438_[12], _0438_[12:11], _0438_[11], _0438_[11], _0438_[11], _0438_[11], _0438_[11], _0438_[11], _0438_[11], _0438_[11], _0438_[11], _0438_[11], _0438_[11], _0438_[11], _0438_[11], _0438_[11], _0438_[11], _0438_[11], _0438_[11], _0438_[11], _0438_[11], _0438_[11:10], _0438_[10], _0438_[10], _0438_[10], _0438_[10], _0438_[10], _0438_[10], _0438_[10], _0438_[10], _0438_[10], _0438_[10], _0438_[10], _0438_[10], _0438_[10], _0438_[10], _0438_[10], _0438_[10], _0438_[10], _0438_[10], _0438_[10], _0438_[10], _0438_[10:9], _0438_[9], _0438_[9], _0438_[9], _0438_[9], _0438_[9], _0438_[9], _0438_[9], _0438_[9], _0438_[9], _0438_[9], _0438_[9], _0438_[9], _0438_[9], _0438_[9], _0438_[9], _0438_[9], _0438_[9], _0438_[9], _0438_[9], _0438_[9], _0438_[9], _0438_[9:8], _0438_[8], _0438_[8], _0438_[8], _0438_[8], _0438_[8], _0438_[8], _0438_[8], _0438_[8], _0438_[8], _0438_[8], _0438_[8], _0438_[8], _0438_[8], _0438_[8], _0438_[8], _0438_[8], _0438_[8], _0438_[8], _0438_[8], _0438_[8], _0438_[8], _0438_[8], _0438_[8:7], _0438_[7], _0438_[7], _0438_[7], _0438_[7], _0438_[7], _0438_[7], _0438_[7], _0438_[7], _0438_[7], _0438_[7], _0438_[7], _0438_[7], _0438_[7], _0438_[7], _0438_[7], _0438_[7], _0438_[7], _0438_[7], _0438_[7], _0438_[7], _0438_[7], _0438_[7], _0438_[7], _0438_[7:6], _0438_[6], _0438_[6], _0438_[6], _0438_[6], _0438_[6], _0438_[6], _0438_[6], _0438_[6], _0438_[6], _0438_[6], _0438_[6], _0438_[6], _0438_[6], _0438_[6], _0438_[6], _0438_[6], _0438_[6], _0438_[6], _0438_[6], _0438_[6], _0438_[6], _0438_[6], _0438_[6], _0438_[6], _0438_[6:5], _0438_[5], _0438_[5], _0438_[5], _0438_[5], _0438_[5], _0438_[5], _0438_[5], _0438_[5], _0438_[5], _0438_[5], _0438_[5], _0438_[5], _0438_[5], _0438_[5], _0438_[5], _0438_[5], _0438_[5], _0438_[5], _0438_[5], _0438_[5], _0438_[5], _0438_[5], _0438_[5], _0438_[5], _0438_[5], _0438_[5:4], _0438_[4], _0438_[4], _0438_[4], _0438_[4], _0438_[4], _0438_[4], _0438_[4], _0438_[4], _0438_[4], _0438_[4], _0438_[4], _0438_[4], _0438_[4], _0438_[4], _0438_[4], _0438_[4], _0438_[4], _0438_[4], _0438_[4], _0438_[4], _0438_[4], _0438_[4], _0438_[4], _0438_[4], _0438_[4], _0438_[4], _0438_[4:3], _0438_[3], _0438_[3], _0438_[3], _0438_[3], _0438_[3], _0438_[3], _0438_[3], _0438_[3], _0438_[3], _0438_[3], _0438_[3], _0438_[3], _0438_[3], _0438_[3], _0438_[3], _0438_[3], _0438_[3], _0438_[3], _0438_[3], _0438_[3], _0438_[3], _0438_[3], _0438_[3], _0438_[3], _0438_[3], _0438_[3], _0438_[3], _0438_[3:2], _0438_[2], _0438_[2], _0438_[2], _0438_[2], _0438_[2], _0438_[2], _0438_[2], _0438_[2], _0438_[2], _0438_[2], _0438_[2], _0438_[2], _0438_[2], _0438_[2], _0438_[2], _0438_[2], _0438_[2], _0438_[2], _0438_[2], _0438_[2], _0438_[2], _0438_[2], _0438_[2], _0438_[2], _0438_[2], _0438_[2], _0438_[2], _0438_[2], _0438_[2:1], _0438_[1], _0438_[1], _0438_[1], _0438_[1], _0438_[1], _0438_[1], _0438_[1], _0438_[1], _0438_[1], _0438_[1], _0438_[1], _0438_[1], _0438_[1], _0438_[1], _0438_[1], _0438_[1], _0438_[1], _0438_[1], _0438_[1], _0438_[1], _0438_[1], _0438_[1], _0438_[1], _0438_[1], _0438_[1], _0438_[1], _0438_[1], _0438_[1], _0438_[1], _0438_[1:0], _0438_[0], _0438_[0], _0438_[0], _0438_[0], _0438_[0], _0438_[0], _0438_[0], _0438_[0], _0438_[0], _0438_[0], _0438_[0], _0438_[0], _0438_[0], _0438_[0], _0438_[0], _0438_[0], _0438_[0], _0438_[0], _0438_[0], _0438_[0], _0438_[0], _0438_[0], _0438_[0], _0438_[0], _0438_[0], _0438_[0], _0438_[0], _0438_[0], _0438_[0], _0438_[0], _0438_[0] } | { _0438_[32], _0438_[32:31], _0438_[32:30], _0438_[32:29], _0438_[32:28], _0438_[32:27], _0438_[32:26], _0438_[32:25], _0438_[32:24], _0438_[32:23], _0438_[32:22], _0438_[32:21], _0438_[32:20], _0438_[32:19], _0438_[32:18], _0438_[32:17], _0438_[32:16], _0438_[32:15], _0438_[32:14], _0438_[32:13], _0438_[32:12], _0438_[32:11], _0438_[32:10], _0438_[32:9], _0438_[32:8], _0438_[32:7], _0438_[32:6], _0438_[32:5], _0438_[32:4], _0438_[32:3], _0438_[32:2], _0438_[32:1] };
  assign _0294_ = _0329_ | _0293_;
  assign _0214_ = _0294_ & { _0359_, _0360_, _0359_, _0361_, _0360_, _0359_, _0362_, _0361_, _0360_, _0359_, _0363_, _0362_, _0361_, _0360_, _0359_, _0364_, _0363_, _0362_, _0361_, _0360_, _0359_, _0365_, _0364_, _0363_, _0362_, _0361_, _0360_, _0359_, _0366_, _0365_, _0364_, _0363_, _0362_, _0361_, _0360_, _0359_, _0367_, _0366_, _0365_, _0364_, _0363_, _0362_, _0361_, _0360_, _0359_, _0368_, _0367_, _0366_, _0365_, _0364_, _0363_, _0362_, _0361_, _0360_, _0359_, _0369_, _0368_, _0367_, _0366_, _0365_, _0364_, _0363_, _0362_, _0361_, _0360_, _0359_, _0370_, _0369_, _0368_, _0367_, _0366_, _0365_, _0364_, _0363_, _0362_, _0361_, _0360_, _0359_, _0371_, _0370_, _0369_, _0368_, _0367_, _0366_, _0365_, _0364_, _0363_, _0362_, _0361_, _0360_, _0359_, _0372_, _0371_, _0370_, _0369_, _0368_, _0367_, _0366_, _0365_, _0364_, _0363_, _0362_, _0361_, _0360_, _0359_, _0373_, _0372_, _0371_, _0370_, _0369_, _0368_, _0367_, _0366_, _0365_, _0364_, _0363_, _0362_, _0361_, _0360_, _0359_, _0374_, _0373_, _0372_, _0371_, _0370_, _0369_, _0368_, _0367_, _0366_, _0365_, _0364_, _0363_, _0362_, _0361_, _0360_, _0359_, _0375_, _0374_, _0373_, _0372_, _0371_, _0370_, _0369_, _0368_, _0367_, _0366_, _0365_, _0364_, _0363_, _0362_, _0361_, _0360_, _0359_, _0376_, _0375_, _0374_, _0373_, _0372_, _0371_, _0370_, _0369_, _0368_, _0367_, _0366_, _0365_, _0364_, _0363_, _0362_, _0361_, _0360_, _0359_, _0377_, _0376_, _0375_, _0374_, _0373_, _0372_, _0371_, _0370_, _0369_, _0368_, _0367_, _0366_, _0365_, _0364_, _0363_, _0362_, _0361_, _0360_, _0359_, _0378_, _0377_, _0376_, _0375_, _0374_, _0373_, _0372_, _0371_, _0370_, _0369_, _0368_, _0367_, _0366_, _0365_, _0364_, _0363_, _0362_, _0361_, _0360_, _0359_, _0379_, _0378_, _0377_, _0376_, _0375_, _0374_, _0373_, _0372_, _0371_, _0370_, _0369_, _0368_, _0367_, _0366_, _0365_, _0364_, _0363_, _0362_, _0361_, _0360_, _0359_, _0380_, _0379_, _0378_, _0377_, _0376_, _0375_, _0374_, _0373_, _0372_, _0371_, _0370_, _0369_, _0368_, _0367_, _0366_, _0365_, _0364_, _0363_, _0362_, _0361_, _0360_, _0359_, _0381_, _0380_, _0379_, _0378_, _0377_, _0376_, _0375_, _0374_, _0373_, _0372_, _0371_, _0370_, _0369_, _0368_, _0367_, _0366_, _0365_, _0364_, _0363_, _0362_, _0361_, _0360_, _0359_, _0382_, _0381_, _0380_, _0379_, _0378_, _0377_, _0376_, _0375_, _0374_, _0373_, _0372_, _0371_, _0370_, _0369_, _0368_, _0367_, _0366_, _0365_, _0364_, _0363_, _0362_, _0361_, _0360_, _0359_, _0383_, _0382_, _0381_, _0380_, _0379_, _0378_, _0377_, _0376_, _0375_, _0374_, _0373_, _0372_, _0371_, _0370_, _0369_, _0368_, _0367_, _0366_, _0365_, _0364_, _0363_, _0362_, _0361_, _0360_, _0359_, _0384_, _0383_, _0382_, _0381_, _0380_, _0379_, _0378_, _0377_, _0376_, _0375_, _0374_, _0373_, _0372_, _0371_, _0370_, _0369_, _0368_, _0367_, _0366_, _0365_, _0364_, _0363_, _0362_, _0361_, _0360_, _0359_, _0385_, _0384_, _0383_, _0382_, _0381_, _0380_, _0379_, _0378_, _0377_, _0376_, _0375_, _0374_, _0373_, _0372_, _0371_, _0370_, _0369_, _0368_, _0367_, _0366_, _0365_, _0364_, _0363_, _0362_, _0361_, _0360_, _0359_, _0386_, _0385_, _0384_, _0383_, _0382_, _0381_, _0380_, _0379_, _0378_, _0377_, _0376_, _0375_, _0374_, _0373_, _0372_, _0371_, _0370_, _0369_, _0368_, _0367_, _0366_, _0365_, _0364_, _0363_, _0362_, _0361_, _0360_, _0359_, _0387_, _0386_, _0385_, _0384_, _0383_, _0382_, _0381_, _0380_, _0379_, _0378_, _0377_, _0376_, _0375_, _0374_, _0373_, _0372_, _0371_, _0370_, _0369_, _0368_, _0367_, _0366_, _0365_, _0364_, _0363_, _0362_, _0361_, _0360_, _0359_, _0388_, _0387_, _0386_, _0385_, _0384_, _0383_, _0382_, _0381_, _0380_, _0379_, _0378_, _0377_, _0376_, _0375_, _0374_, _0373_, _0372_, _0371_, _0370_, _0369_, _0368_, _0367_, _0366_, _0365_, _0364_, _0363_, _0362_, _0361_, _0360_, _0359_, _0389_, _0388_, _0387_, _0386_, _0385_, _0384_, _0383_, _0382_, _0381_, _0380_, _0379_, _0378_, _0377_, _0376_, _0375_, _0374_, _0373_, _0372_, _0371_, _0370_, _0369_, _0368_, _0367_, _0366_, _0365_, _0364_, _0363_, _0362_, _0361_, _0360_, _0359_, 1'h0, _0389_, _0388_, _0387_, _0386_, _0385_, _0384_, _0383_, _0382_, _0381_, _0380_, _0379_, _0378_, _0377_, _0376_, _0375_, _0374_, _0373_, _0372_, _0371_, _0370_, _0369_, _0368_, _0367_, _0366_, _0365_, _0364_, _0363_, _0362_, _0361_, _0360_, _0359_ };
  assign _0390_ = { 1'h0, shift_amt_t0[4:0] } >= 32'd33;
  assign _0391_ = { 1'h0, shift_amt_t0[4:0] } >= 32'd32;
  assign _0392_ = { 1'h0, shift_amt_t0[4:0] } >= 32'd31;
  assign _0393_ = { 1'h0, shift_amt_t0[4:0] } >= 32'd30;
  assign _0394_ = { 1'h0, shift_amt_t0[4:0] } >= 32'd29;
  assign _0395_ = { 1'h0, shift_amt_t0[4:0] } >= 32'd28;
  assign _0396_ = { 1'h0, shift_amt_t0[4:0] } >= 32'd27;
  assign _0397_ = { 1'h0, shift_amt_t0[4:0] } >= 32'd26;
  assign _0398_ = { 1'h0, shift_amt_t0[4:0] } >= 32'd25;
  assign _0399_ = { 1'h0, shift_amt_t0[4:0] } >= 32'd24;
  assign _0400_ = { 1'h0, shift_amt_t0[4:0] } >= 32'd23;
  assign _0401_ = { 1'h0, shift_amt_t0[4:0] } >= 32'd22;
  assign _0402_ = { 1'h0, shift_amt_t0[4:0] } >= 32'd21;
  assign _0403_ = { 1'h0, shift_amt_t0[4:0] } >= 32'd20;
  assign _0404_ = { 1'h0, shift_amt_t0[4:0] } >= 32'd19;
  assign _0405_ = { 1'h0, shift_amt_t0[4:0] } >= 32'd18;
  assign _0406_ = { 1'h0, shift_amt_t0[4:0] } >= 32'd17;
  assign _0407_ = { 1'h0, shift_amt_t0[4:0] } >= 32'd16;
  assign _0408_ = { 1'h0, shift_amt_t0[4:0] } >= 32'd15;
  assign _0409_ = { 1'h0, shift_amt_t0[4:0] } >= 32'd14;
  assign _0410_ = { 1'h0, shift_amt_t0[4:0] } >= 32'd13;
  assign _0411_ = { 1'h0, shift_amt_t0[4:0] } >= 32'd12;
  assign _0412_ = { 1'h0, shift_amt_t0[4:0] } >= 32'd11;
  assign _0413_ = { 1'h0, shift_amt_t0[4:0] } >= 32'd10;
  assign _0414_ = { 1'h0, shift_amt_t0[4:0] } >= 32'd9;
  assign _0415_ = { 1'h0, shift_amt_t0[4:0] } >= 32'd8;
  assign _0416_ = { 1'h0, shift_amt_t0[4:0] } >= 32'd7;
  assign _0417_ = { 1'h0, shift_amt_t0[4:0] } >= 32'd6;
  assign _0418_ = { 1'h0, shift_amt_t0[4:0] } >= 32'd5;
  assign _0419_ = { 1'h0, shift_amt_t0[4:0] } >= 32'd4;
  assign _0420_ = { 1'h0, shift_amt_t0[4:0] } >= 32'd3;
  assign _0421_ = { 1'h0, shift_amt_t0[4:0] } >= 32'd2;
  assign _0422_ = { 1'h0, shift_amt_t0[4:0] } >= 32'd1;
  assign _0330_ = _0437_ ^ { _0437_[32], _0437_[32], _0437_[32], _0437_[32], _0437_[32], _0437_[32], _0437_[32], _0437_[32], _0437_[32], _0437_[32], _0437_[32], _0437_[32], _0437_[32], _0437_[32], _0437_[32], _0437_[32], _0437_[32], _0437_[32], _0437_[32], _0437_[32], _0437_[32], _0437_[32], _0437_[32], _0437_[32], _0437_[32], _0437_[32], _0437_[32], _0437_[32], _0437_[32], _0437_[32], _0437_[32], _0437_[32], _0437_[32] };
  assign _0295_ = _0438_ | _0330_;
  assign _0215_ = _0295_ & { _0422_, _0421_, _0420_, _0419_, _0418_, _0417_, _0416_, _0415_, _0414_, _0413_, _0412_, _0411_, _0410_, _0409_, _0408_, _0407_, _0406_, _0405_, _0404_, _0403_, _0402_, _0401_, _0400_, _0399_, _0398_, _0397_, _0396_, _0395_, _0394_, _0393_, _0392_, _0391_, _0390_ };
  assign shift_result_ext_t0[0] = | { _0215_[0], _0214_[31:0], _0438_[0] };
  assign shift_result_ext_t0[1] = | { _0215_[1], _0214_[62:32], _0438_[1] };
  assign shift_result_ext_t0[2] = | { _0215_[2], _0214_[92:63], _0438_[2] };
  assign shift_result_ext_t0[3] = | { _0215_[3], _0214_[121:93], _0438_[3] };
  assign shift_result_ext_t0[4] = | { _0215_[4], _0214_[149:122], _0438_[4] };
  assign shift_result_ext_t0[5] = | { _0215_[5], _0214_[176:150], _0438_[5] };
  assign shift_result_ext_t0[6] = | { _0215_[6], _0214_[202:177], _0438_[6] };
  assign shift_result_ext_t0[7] = | { _0215_[7], _0214_[227:203], _0438_[7] };
  assign shift_result_ext_t0[8] = | { _0215_[8], _0214_[251:228], _0438_[8] };
  assign shift_result_ext_t0[9] = | { _0215_[9], _0214_[274:252], _0438_[9] };
  assign shift_result_ext_t0[10] = | { _0215_[10], _0214_[296:275], _0438_[10] };
  assign shift_result_ext_t0[11] = | { _0215_[11], _0214_[317:297], _0438_[11] };
  assign shift_result_ext_t0[12] = | { _0215_[12], _0214_[337:318], _0438_[12] };
  assign shift_result_ext_t0[13] = | { _0215_[13], _0214_[356:338], _0438_[13] };
  assign shift_result_ext_t0[14] = | { _0215_[14], _0214_[374:357], _0438_[14] };
  assign shift_result_ext_t0[15] = | { _0215_[15], _0214_[391:375], _0438_[15] };
  assign shift_result_ext_t0[16] = | { _0215_[16], _0214_[407:392], _0438_[16] };
  assign shift_result_ext_t0[17] = | { _0215_[17], _0214_[422:408], _0438_[17] };
  assign shift_result_ext_t0[18] = | { _0215_[18], _0214_[436:423], _0438_[18] };
  assign shift_result_ext_t0[19] = | { _0215_[19], _0214_[449:437], _0438_[19] };
  assign shift_result_ext_t0[20] = | { _0215_[20], _0214_[461:450], _0438_[20] };
  assign shift_result_ext_t0[21] = | { _0215_[21], _0214_[472:462], _0438_[21] };
  assign shift_result_ext_t0[22] = | { _0215_[22], _0214_[482:473], _0438_[22] };
  assign shift_result_ext_t0[23] = | { _0215_[23], _0214_[491:483], _0438_[23] };
  assign shift_result_ext_t0[24] = | { _0215_[24], _0214_[499:492], _0438_[24] };
  assign shift_result_ext_t0[25] = | { _0215_[25], _0214_[506:500], _0438_[25] };
  assign shift_result_ext_t0[26] = | { _0215_[26], _0214_[512:507], _0438_[26] };
  assign shift_result_ext_t0[27] = | { _0215_[27], _0214_[517:513], _0438_[27] };
  assign shift_result_ext_t0[28] = | { _0215_[28], _0214_[521:518], _0438_[28] };
  assign shift_result_ext_t0[29] = | { _0215_[29], _0214_[524:522], _0438_[29] };
  assign shift_result_ext_t0[30] = | { _0215_[30], _0214_[526:525], _0438_[30] };
  assign shift_result_ext_t0[31] = | { _0215_[31], _0214_[527], _0438_[31] };
  assign _0039_ = ~ { 1'h0, shift_amt_t0[4:0] };
  assign _0182_ = { 1'h0, shift_amt[4:0] } & _0039_;
  assign _0437_ = $signed({ _0000_, shift_operand }) >>> _0182_;
  assign _0438_ = $signed({ _0001_, shift_operand_t0 }) >>> _0182_;
  assign _0040_ = ~ { 27'h0000000, operand_b_i_t0[4:0] };
  assign _0216_ = { 27'h0000000, operand_b_i[4:0] } & _0040_;
  assign _0296_ = { 27'h0000000, operand_b_i[4:0] } | { 27'h0000000, operand_b_i_t0[4:0] };
  assign _0425_ = 32'd32 - _0216_;
  assign _0426_ = 32'd32 - _0296_;
  assign _0297_ = _0425_ ^ _0426_;
  assign { _0501_[31:6], shift_amt_compl_t0 } = _0297_ | { 27'h0000000, operand_b_i_t0[4:0] };
  assign bwlogic_xor_result_t0 = operand_a_i_t0 | operand_b_i_t0;
  assign _0503_ = operand_a_i_t0[31] | operand_b_i_t0[31];
  assign _0505_ = operand_a_i_t0[31] | cmp_signed_t0;
  assign is_equal_result_o = ! adder_result_ext_o[32:1];
  assign _0447_ = ~ adder_result_ext_o[32];
  assign adder_op_b_negate = operator_i[5] ? _0450_ : _0448_;
  assign _0448_ = operator_i[4] ? _0454_ : _0452_;
  assign _0450_ = operator_i[4] ? 1'h0 : _0315_;
  assign _0452_ = operator_i[3] ? 1'h0 : _0316_;
  assign _0454_ = operator_i[3] ? _0460_ : _0458_;
  assign _0315_ = operator_i[3] ? 1'h0 : _0318_;
  assign _0316_ = operator_i[2] ? 1'h0 : _0319_;
  assign _0458_ = operator_i[2] ? 1'h1 : _0464_;
  assign _0460_ = operator_i[2] ? _0466_ : 1'h1;
  assign _0318_ = operator_i[2] ? _0320_ : 1'h0;
  assign _0319_ = operator_i[1] ? 1'h0 : _0321_;
  assign _0464_ = operator_i[1] ? _0321_ : 1'h0;
  assign _0466_ = operator_i[1] ? 1'h0 : _0322_;
  assign _0320_ = operator_i[1] ? _0322_ : _0321_;
  assign _0321_ = operator_i[0] ? 1'h1 : 1'h0;
  assign _0322_ = operator_i[0] ? 1'h0 : 1'h1;
  assign _0469_ = ~ is_equal_result_o;
  assign _0470_ = ~ is_greater_equal;
  assign bwlogic_or_result = operand_a_i | operand_b_i;
  assign bwlogic_or = _0439_ | _0441_;
  assign bwlogic_and = _0443_ | _0445_;
  assign _0473_ = | _0471_;
  assign _0471_[0] = operator_i == 6'h17;
  assign _0477_ = | { _0475_[4:3], _0475_[1:0], shift_arith };
  assign _0475_[1] = operator_i == 6'h09;
  assign shift_arith = operator_i == 6'h08;
  assign _0475_[3] = operator_i == 6'h0c;
  assign _0475_[4] = operator_i == 6'h0b;
  assign _0481_ = | _0479_;
  assign _0479_[0] = ! operator_i;
  assign _0479_[1] = operator_i == 6'h01;
  assign _0485_ = | { _0483_[1:0], _0445_, _0443_, _0441_, _0439_ };
  assign _0483_[0] = operator_i == 6'h02;
  assign _0483_[1] = operator_i == 6'h05;
  assign _0439_ = operator_i == 6'h03;
  assign _0441_ = operator_i == 6'h06;
  assign _0443_ = operator_i == 6'h04;
  assign _0445_ = operator_i == 6'h07;
  assign _0487_ = bwlogic_and ? bwlogic_and_result : bwlogic_xor_result;
  assign bwlogic_result = bwlogic_or ? bwlogic_or_result : _0487_;
  assign shift_left = _0475_[0] ? 1'h1 : 1'h0;
  assign _0475_[0] = operator_i == 6'h0a;
  assign _0491_ = | { _0489_[3:2], _0471_[7:4] };
  assign _0471_[4] = operator_i == 6'h13;
  assign _0471_[5] = operator_i == 6'h14;
  assign _0489_[2] = operator_i == 6'h19;
  assign _0489_[3] = operator_i == 6'h1a;
  assign _0471_[6] = operator_i == 6'h25;
  assign _0471_[7] = operator_i == 6'h26;
  assign _0495_ = | { _0493_[3:2], _0471_[3:2] };
  assign _0471_[2] = operator_i == 6'h15;
  assign _0471_[3] = operator_i == 6'h16;
  assign _0493_[2] = operator_i == 6'h1b;
  assign _0493_[3] = operator_i == 6'h1c;
  assign _0471_[1] = operator_i == 6'h18;
  assign is_greater_equal = _0502_ ? _0504_ : _0447_;
  assign cmp_signed = _0497_ ? 1'h1 : 1'h0;
  assign _0497_ = | { _0493_[2], _0489_[2], _0471_[6], _0471_[4], _0471_[2] };
  assign _0498_ = adder_op_b_negate ? operand_b_neg : { operand_b_i, 1'h0 };
  assign adder_in_b = multdiv_sel_i ? multdiv_operand_b_i : _0498_;
  assign shift_result_ext = $signed({ _0000_, shift_operand }) >>> shift_amt[4:0];
  assign { _0500_[31:6], shift_amt_compl } = 32'd32 - operand_b_i[4:0];
  assign shift_amt[4:0] = instr_first_cycle_i ? operand_b_i[4:0] : shift_amt_compl[4:0];
  assign shift_operand = shift_left ? { operand_a_i[0], operand_a_i[1], operand_a_i[2], operand_a_i[3], operand_a_i[4], operand_a_i[5], operand_a_i[6], operand_a_i[7], operand_a_i[8], operand_a_i[9], operand_a_i[10], operand_a_i[11], operand_a_i[12], operand_a_i[13], operand_a_i[14], operand_a_i[15], operand_a_i[16], operand_a_i[17], operand_a_i[18], operand_a_i[19], operand_a_i[20], operand_a_i[21], operand_a_i[22], operand_a_i[23], operand_a_i[24], operand_a_i[25], operand_a_i[26], operand_a_i[27], operand_a_i[28], operand_a_i[29], operand_a_i[30], operand_a_i[31] } : operand_a_i;
  assign shift_result = shift_left ? { shift_result_ext[0], shift_result_ext[1], shift_result_ext[2], shift_result_ext[3], shift_result_ext[4], shift_result_ext[5], shift_result_ext[6], shift_result_ext[7], shift_result_ext[8], shift_result_ext[9], shift_result_ext[10], shift_result_ext[11], shift_result_ext[12], shift_result_ext[13], shift_result_ext[14], shift_result_ext[15], shift_result_ext[16], shift_result_ext[17], shift_result_ext[18], shift_result_ext[19], shift_result_ext[20], shift_result_ext[21], shift_result_ext[22], shift_result_ext[23], shift_result_ext[24], shift_result_ext[25], shift_result_ext[26], shift_result_ext[27], shift_result_ext[28], shift_result_ext[29], shift_result_ext[30], shift_result_ext[31] } : shift_result_ext[31:0];
  assign adder_in_a = multdiv_sel_i ? multdiv_operand_a_i : { operand_a_i, 1'h1 };
  assign bwlogic_xor_result = operand_a_i ^ operand_b_i;
  assign operand_b_neg = { operand_b_i, 1'h0 } ^ 33'h1ffffffff;
  assign _0502_ = operand_a_i[31] ^ operand_b_i[31];
  assign _0504_ = operand_a_i[31] ^ cmp_signed;
  assign _0475_[2] = shift_arith;
  assign { _0476_[2], _0476_[0] } = { shift_arith_t0, shift_left_t0 };
  assign _0483_[5:2] = { _0445_, _0443_, _0441_, _0439_ };
  assign _0484_[5:2] = { _0446_, _0444_, _0442_, _0440_ };
  assign { _0489_[5:4], _0489_[1:0] } = _0471_[7:4];
  assign { _0490_[5:4], _0490_[1:0] } = _0472_[7:4];
  assign _0493_[1:0] = _0471_[3:2];
  assign _0494_[1:0] = _0472_[3:2];
  assign _0500_[5:0] = shift_amt_compl;
  assign _0501_[5:0] = shift_amt_compl_t0;
  assign adder_result_o = adder_result_ext_o[32:1];
  assign adder_result_o_t0 = adder_result_ext_o_t0[32:1];
  assign imd_val_d_o = 64'h0000000000000000;
  assign imd_val_d_o_t0 = 64'h0000000000000000;
  assign imd_val_we_o = 2'h0;
  assign imd_val_we_o_t0 = 2'h0;
  assign shift_amt[5] = 1'h0;
  assign shift_amt_t0[5] = 1'h0;
endmodule






module paramodauxy_ibex_controllerWritebackStage11BranchPredictor10 (clk_i, rst_ni, ctrl_busy_o, illegal_insn_i, ecall_insn_i, mret_insn_i, dret_insn_i, wfi_insn_i, ebrk_insn_i, csr_pipe_flush_i, instr_valid_i, instr_i, instr_compressed_i, instr_is_compressed_i, instr_bp_taken_i, instr_fetch_err_i, instr_fetch_err_plus2_i, pc_id_i, instr_valid_clear_o, id_in_ready_o, controller_run_o
, instr_req_o, pc_set_o, pc_set_spec_o, pc_mux_o, nt_branch_mispredict_o, exc_pc_mux_o, exc_cause_o, lsu_addr_last_i, load_err_i, store_err_i, wb_exception_o, branch_set_i, branch_set_spec_i, branch_not_set_i, jump_set_i, csr_mstatus_mie_i, irq_pending_i, irqs_i, irq_nm_i, nmi_mode_o, debug_req_i
, debug_cause_o, debug_csr_save_o, debug_mode_o, debug_single_step_i, debug_ebreakm_i, debug_ebreaku_i, trigger_match_i, csr_save_if_o, csr_save_id_o, csr_save_wb_o, csr_restore_mret_id_o, csr_restore_dret_id_o, csr_save_cause_o, csr_mtval_o, priv_mode_i, csr_mstatus_tw_i, stall_id_i, stall_wb_i, flush_id_o, ready_wb_i, perf_jump_o
, perf_tbranch_o, instr_req_o_t0, instr_i_t0, branch_not_set_i_t0, branch_set_i_t0, branch_set_spec_i_t0, controller_run_o_t0, csr_mstatus_mie_i_t0, csr_mstatus_tw_i_t0, csr_mtval_o_t0, csr_pipe_flush_i_t0, csr_restore_dret_id_o_t0, csr_restore_mret_id_o_t0, csr_save_cause_o_t0, csr_save_id_o_t0, csr_save_if_o_t0, csr_save_wb_o_t0, ctrl_busy_o_t0, debug_cause_o_t0, debug_csr_save_o_t0, debug_ebreakm_i_t0
, debug_ebreaku_i_t0, debug_mode_o_t0, debug_req_i_t0, debug_single_step_i_t0, dret_insn_i_t0, ebrk_insn_i_t0, ecall_insn_i_t0, exc_cause_o_t0, exc_pc_mux_o_t0, flush_id_o_t0, id_in_ready_o_t0, illegal_insn_i_t0, instr_bp_taken_i_t0, instr_compressed_i_t0, instr_fetch_err_i_t0, instr_fetch_err_plus2_i_t0, instr_is_compressed_i_t0, instr_valid_clear_o_t0, instr_valid_i_t0, irq_nm_i_t0, irq_pending_i_t0
, irqs_i_t0, jump_set_i_t0, load_err_i_t0, lsu_addr_last_i_t0, mret_insn_i_t0, nmi_mode_o_t0, nt_branch_mispredict_o_t0, pc_id_i_t0, pc_mux_o_t0, pc_set_o_t0, pc_set_spec_o_t0, perf_jump_o_t0, perf_tbranch_o_t0, priv_mode_i_t0, ready_wb_i_t0, stall_id_i_t0, stall_wb_i_t0, store_err_i_t0, trigger_match_i_t0, wb_exception_o_t0, wfi_insn_i_t0
);
  wire [3:0] _0000_;
  wire [3:0] _0001_;
  wire [3:0] _0002_;
  wire [3:0] _0003_;
  wire [3:0] _0004_;
  wire [3:0] _0005_;
  wire [3:0] _0006_;
  wire [3:0] _0007_;
  wire [3:0] _0008_;
  wire [3:0] _0009_;
  wire [3:0] _0010_;
  wire [3:0] _0011_;
  wire [3:0] _0012_;
  wire [3:0] _0013_;
  wire [3:0] _0014_;
  wire [3:0] _0015_;
  wire [3:0] _0016_;
  wire [3:0] _0017_;
  wire [3:0] _0018_;
  wire [3:0] _0019_;
  wire [3:0] _0020_;
  wire [3:0] _0021_;
  wire [3:0] _0022_;
  wire [3:0] _0023_;
  wire [3:0] _0024_;
  wire [3:0] _0025_;
  wire [3:0] _0026_;
  wire [3:0] _0027_;
  wire [31:0] _0028_;
  wire [31:0] _0029_;
  wire _0030_;
  wire _0031_;
  wire _0032_;
  wire _0033_;
  wire _0034_;
  wire _0035_;
  wire _0036_;
  wire _0037_;
  wire _0038_;
  wire _0039_;
  wire _0040_;
  wire [3:0] _0041_;
  wire [3:0] _0042_;
  wire [2:0] _0043_;
  wire [2:0] _0044_;
  wire _0045_;
  wire _0046_;
  wire _0047_;
  wire _0048_;
  wire _0049_;
  wire [5:0] _0050_;
  wire [5:0] _0051_;
  wire [1:0] _0052_;
  wire [1:0] _0053_;
  wire _0054_;
  wire _0055_;
  wire _0056_;
  wire _0057_;
  wire _0058_;
  wire _0059_;
  wire _0060_;
  wire [3:0] _0061_;
  wire [3:0] _0062_;
  wire _0063_;
  wire [2:0] _0064_;
  wire [2:0] _0065_;
  wire _0066_;
  wire _0067_;
  wire _0068_;
  wire _0069_;
  wire _0070_;
  wire _0071_;
  wire _0072_;
  wire _0073_;
  wire _0074_;
  wire [31:0] _0075_;
  wire [31:0] _0076_;
  wire _0077_;
  wire _0078_;
  wire _0079_;
  wire _0080_;
  wire _0081_;
  wire _0082_;
  wire _0083_;
  wire [3:0] _0084_;
  wire [3:0] _0085_;
  wire [2:0] _0086_;
  wire [2:0] _0087_;
  wire _0088_;
  wire _0089_;
  wire _0090_;
  wire _0091_;
  wire _0092_;
  wire [5:0] _0093_;
  wire [5:0] _0094_;
  wire _0095_;
  wire _0096_;
  wire _0097_;
  wire _0098_;
  wire _0099_;
  wire _0100_;
  wire _0101_;
  wire [3:0] _0102_;
  wire [3:0] _0103_;
  wire _0104_;
  wire [2:0] _0105_;
  wire [2:0] _0106_;
  wire _0107_;
  wire _0108_;
  wire _0109_;
  wire _0110_;
  wire [3:0] _0111_;
  wire [3:0] _0112_;
  wire _0113_;
  wire _0114_;
  wire _0115_;
  wire _0116_;
  wire _0117_;
  wire [5:0] _0118_;
  wire [5:0] _0119_;
  wire _0120_;
  wire _0121_;
  wire _0122_;
  wire _0123_;
  wire _0124_;
  wire [3:0] _0125_;
  wire [3:0] _0126_;
  wire _0127_;
  wire [2:0] _0128_;
  wire [2:0] _0129_;
  wire _0130_;
  wire _0131_;
  wire _0132_;
  wire _0133_;
  wire [3:0] _0134_;
  wire [3:0] _0135_;
  wire _0136_;
  wire _0137_;
  wire _0138_;
  wire [5:0] _0139_;
  wire [5:0] _0140_;
  wire _0141_;
  wire _0142_;
  wire [3:0] _0143_;
  wire [3:0] _0144_;
  wire _0145_;
  wire _0146_;
  wire _0147_;
  wire [3:0] _0148_;
  wire [3:0] _0149_;
  wire _0150_;
  wire [5:0] _0151_;
  wire [5:0] _0152_;
  wire _0153_;
  wire _0154_;
  wire [3:0] _0155_;
  wire [3:0] _0156_;
  wire [3:0] _0157_;
  wire [3:0] _0158_;
  wire [5:0] _0159_;
  wire [5:0] _0160_;
  wire _0161_;
  wire _0162_;
  wire [3:0] _0163_;
  wire [3:0] _0164_;
  wire _0165_;
  wire _0166_;
  wire [3:0] _0167_;
  wire [3:0] _0168_;
  wire [5:0] _0169_;
  wire [5:0] _0170_;
  wire [3:0] _0171_;
  wire [3:0] _0172_;
  wire [3:0] _0173_;
  wire [3:0] _0174_;
  wire [5:0] _0175_;
  wire [5:0] _0176_;
  wire [3:0] _0177_;
  wire [3:0] _0178_;
  wire [31:0] _0179_;
  wire [31:0] _0180_;
  wire _0181_;
  wire _0182_;
  wire _0183_;
  wire _0184_;
  wire _0185_;
  wire _0186_;
  wire _0187_;
  wire _0188_;
  wire _0189_;
  wire _0190_;
  wire _0191_;
  wire _0192_;
  wire _0193_;
  wire _0194_;
  wire _0195_;
  wire _0196_;
  wire _0197_;
  wire _0198_;
  wire _0199_;
  wire _0200_;
  wire _0201_;
  wire _0202_;
  wire _0203_;
  wire _0204_;
  wire _0205_;
  wire _0206_;
  wire _0207_;
  wire _0208_;
  wire _0209_;
  wire _0210_;
  wire _0211_;
  wire _0212_;
  wire _0213_;
  wire _0214_;
  wire _0215_;
  wire _0216_;
  wire _0217_;
  wire _0218_;
  wire _0219_;
  wire _0220_;
  wire _0221_;
  wire _0222_;
  wire _0223_;
  wire _0224_;
  wire _0225_;
  wire _0226_;
  wire _0227_;
  wire _0228_;
  wire _0229_;
  wire [31:0] _0230_;
  wire _0231_;
  wire _0232_;
  wire _0233_;
  wire [3:0] _0234_;
  wire [2:0] _0235_;
  wire [1:0] _0236_;
  wire [1:0] _0237_;
  wire [1:0] _0238_;
  wire [2:0] _0239_;
  wire [1:0] _0240_;
  wire [3:0] _0241_;
  wire [1:0] _0242_;
  wire [3:0] _0243_;
  wire [3:0] _0244_;
  wire [6:0] _0245_;
  wire [2:0] _0246_;
  wire [2:0] _0247_;
  wire [1:0] _0248_;
  wire _0249_;
  wire _0250_;
  wire _0251_;
  wire _0252_;
  wire _0253_;
  wire _0254_;
  wire _0255_;
  wire _0256_;
  wire [2:0] _0257_;
  wire [3:0] _0258_;
  wire [3:0] _0259_;
  wire [3:0] _0260_;
  wire [3:0] _0261_;
  wire [3:0] _0262_;
  wire [3:0] _0263_;
  wire [3:0] _0264_;
  wire [3:0] _0265_;
  wire _0266_;
  wire _0267_;
  wire [2:0] _0268_;
  wire [2:0] _0269_;
  wire [2:0] _0270_;
  wire _0271_;
  wire _0272_;
  wire _0273_;
  wire [5:0] _0274_;
  wire [5:0] _0275_;
  wire [1:0] _0276_;
  wire [1:0] _0277_;
  wire [1:0] _0278_;
  wire _0279_;
  wire _0280_;
  wire _0281_;
  wire _0282_;
  wire _0283_;
  wire _0284_;
  wire _0285_;
  wire _0286_;
  wire _0287_;
  wire _0288_;
  wire _0289_;
  wire _0290_;
  wire _0291_;
  wire _0292_;
  wire _0293_;
  wire _0294_;
  wire _0295_;
  wire _0296_;
  wire _0297_;
  wire [3:0] _0298_;
  wire [14:0] _0299_;
  wire _0300_;
  wire _0301_;
  wire _0302_;
  wire _0303_;
  wire _0304_;
  wire _0305_;
  wire _0306_;
  wire _0307_;
  wire _0308_;
  wire _0309_;
  wire _0310_;
  wire _0311_;
  wire _0312_;
  wire _0313_;
  wire _0314_;
  wire _0315_;
  wire _0316_;
  wire _0317_;
  wire _0318_;
  wire _0319_;
  wire _0320_;
  wire _0321_;
  wire _0322_;
  wire _0323_;
  wire _0324_;
  wire _0325_;
  wire _0326_;
  wire _0327_;
  wire _0328_;
  wire _0329_;
  wire _0330_;
  wire _0331_;
  wire _0332_;
  wire _0333_;
  wire _0334_;
  wire _0335_;
  wire _0336_;
  wire _0337_;
  wire [3:0] _0338_;
  wire [3:0] _0339_;
  wire [3:0] _0340_;
  wire [2:0] _0341_;
  wire [3:0] _0342_;
  wire [2:0] _0343_;
  wire [3:0] _0344_;
  wire [3:0] _0345_;
  wire _0346_;
  wire [5:0] _0347_;
  wire [31:0] _0348_;
  wire [31:0] _0349_;
  wire [31:0] _0350_;
  wire [31:0] _0351_;
  wire [31:0] _0352_;
  wire [31:0] _0353_;
  wire [5:0] _0354_;
  wire [5:0] _0355_;
  wire [5:0] _0356_;
  wire [5:0] _0357_;
  wire [5:0] _0358_;
  wire [5:0] _0359_;
  wire [3:0] _0360_;
  wire [3:0] _0361_;
  wire [3:0] _0362_;
  wire [3:0] _0363_;
  wire _0364_;
  wire _0365_;
  wire _0366_;
  wire _0367_;
  wire [3:0] _0368_;
  wire _0369_;
  wire [31:0] _0370_;
  wire [5:0] _0371_;
  wire [1:0] _0372_;
  wire [2:0] _0373_;
  wire [2:0] _0374_;
  wire [2:0] _0375_;
  wire [5:0] _0376_;
  wire [5:0] _0377_;
  wire [5:0] _0378_;
  wire [5:0] _0379_;
  wire [5:0] _0380_;
  wire [3:0] _0381_;
  wire [3:0] _0382_;
  wire _0383_;
  wire [3:0] _0384_;
  wire [3:0] _0385_;
  wire [3:0] _0386_;
  wire [3:0] _0387_;
  wire [3:0] _0388_;
  wire [2:0] _0389_;
  wire [31:0] _0390_;
  wire [3:0] _0391_;
  wire [3:0] _0392_;
  wire [3:0] _0393_;
  wire [3:0] _0394_;
  wire [3:0] _0395_;
  wire [3:0] _0396_;
  wire [3:0] _0397_;
  wire [3:0] _0398_;
  wire [3:0] _0399_;
  wire [3:0] _0400_;
  wire [3:0] _0401_;
  wire [3:0] _0402_;
  wire [3:0] _0403_;
  wire [3:0] _0404_;
  wire _0405_;
  wire [1:0] _0406_;
  wire [31:0] _0407_;
  wire [31:0] _0408_;
  wire [5:0] _0409_;
  wire _0410_;
  wire _0411_;
  wire _0412_;
  wire _0413_;
  wire _0414_;
  wire _0415_;
  wire _0416_;
  wire _0417_;
  wire _0418_;
  wire _0419_;
  wire _0420_;
  wire _0421_;
  wire _0422_;
  wire _0423_;
  wire _0424_;
  wire _0425_;
  wire _0426_;
  wire _0427_;
  wire _0428_;
  wire _0429_;
  wire _0430_;
  wire _0431_;
  wire _0432_;
  wire _0433_;
  wire _0434_;
  wire _0435_;
  wire _0436_;
  wire _0437_;
  wire _0438_;
  wire _0439_;
  wire _0440_;
  wire _0441_;
  wire _0442_;
  wire _0443_;
  wire _0444_;
  wire _0445_;
  wire _0446_;
  wire _0447_;
  wire _0448_;
  wire _0449_;
  wire _0450_;
  wire _0451_;
  wire _0452_;
  wire _0453_;
  wire _0454_;
  wire _0455_;
  wire _0456_;
  wire _0457_;
  wire _0458_;
  wire _0459_;
  wire _0460_;
  wire _0461_;
  wire [31:0] _0462_;
  wire _0463_;
  wire _0464_;
  wire _0465_;
  wire _0466_;
  wire _0467_;
  wire _0468_;
  wire _0469_;
  wire _0470_;
  wire _0471_;
  wire _0472_;
  wire _0473_;
  wire _0474_;
  wire _0475_;
  wire _0476_;
  wire _0477_;
  wire _0478_;
  wire _0479_;
  wire _0480_;
  wire _0481_;
  wire _0482_;
  wire _0483_;
  wire _0484_;
  wire _0485_;
  wire _0486_;
  wire _0487_;
  wire _0488_;
  wire _0489_;
  wire _0490_;
  wire _0491_;
  wire _0492_;
  wire _0493_;
  wire _0494_;
  wire _0495_;
  wire _0496_;
  wire _0497_;
  wire _0498_;
  wire _0499_;
  wire _0500_;
  wire _0501_;
  wire _0502_;
  wire _0503_;
  wire _0504_;
  wire _0505_;
  wire _0506_;
  wire _0507_;
  wire _0508_;
  wire _0509_;
  wire _0510_;
  wire _0511_;
  wire _0512_;
  wire _0513_;
  wire _0514_;
  wire _0515_;
  wire _0516_;
  wire _0517_;
  wire _0518_;
  wire _0519_;
  wire _0520_;
  wire _0521_;
  wire _0522_;
  wire _0523_;
  wire _0524_;
  wire _0525_;
  wire _0526_;
  wire _0527_;
  wire _0528_;
  wire [3:0] _0529_;
  wire [3:0] _0530_;
  wire [3:0] _0531_;
  wire [3:0] _0532_;
  wire [3:0] _0533_;
  wire [2:0] _0534_;
  wire [2:0] _0535_;
  wire [1:0] _0536_;
  wire [1:0] _0537_;
  wire [1:0] _0538_;
  wire [2:0] _0539_;
  wire [1:0] _0540_;
  wire [1:0] _0541_;
  wire [2:0] _0542_;
  wire [2:0] _0543_;
  wire [1:0] _0544_;
  wire [3:0] _0545_;
  wire [3:0] _0546_;
  wire [1:0] _0547_;
  wire [1:0] _0548_;
  wire [3:0] _0549_;
  wire [3:0] _0550_;
  wire [6:0] _0551_;
  wire [2:0] _0552_;
  wire [2:0] _0553_;
  wire [1:0] _0554_;
  wire _0555_;
  wire _0556_;
  wire _0557_;
  wire _0558_;
  wire _0559_;
  wire _0560_;
  wire _0561_;
  wire _0562_;
  wire _0563_;
  wire _0564_;
  wire _0565_;
  wire _0566_;
  wire _0567_;
  wire _0568_;
  wire _0569_;
  wire [2:0] _0570_;
  wire [3:0] _0571_;
  wire [3:0] _0572_;
  wire [3:0] _0573_;
  wire [3:0] _0574_;
  wire [3:0] _0575_;
  wire [3:0] _0576_;
  wire [3:0] _0577_;
  wire [3:0] _0578_;
  wire [3:0] _0579_;
  wire [3:0] _0580_;
  wire [3:0] _0581_;
  wire [3:0] _0582_;
  wire [3:0] _0583_;
  wire [3:0] _0584_;
  wire [3:0] _0585_;
  wire [3:0] _0586_;
  wire [3:0] _0587_;
  wire [3:0] _0588_;
  wire [3:0] _0589_;
  wire [3:0] _0590_;
  wire [3:0] _0591_;
  wire [3:0] _0592_;
  wire [3:0] _0593_;
  wire [3:0] _0594_;
  wire _0595_;
  wire _0596_;
  wire _0597_;
  wire _0598_;
  wire _0599_;
  wire _0600_;
  wire _0601_;
  wire _0602_;
  wire _0603_;
  wire _0604_;
  wire _0605_;
  wire _0606_;
  wire _0607_;
  wire _0608_;
  wire _0609_;
  wire _0610_;
  wire [2:0] _0611_;
  wire [2:0] _0612_;
  wire [2:0] _0613_;
  wire [2:0] _0614_;
  wire [2:0] _0615_;
  wire [2:0] _0616_;
  wire [2:0] _0617_;
  wire [2:0] _0618_;
  wire [2:0] _0619_;
  wire _0620_;
  wire _0621_;
  wire _0622_;
  wire _0623_;
  wire _0624_;
  wire _0625_;
  wire _0626_;
  wire _0627_;
  wire _0628_;
  wire _0629_;
  wire _0630_;
  wire _0631_;
  wire _0632_;
  wire _0633_;
  wire _0634_;
  wire _0635_;
  wire _0636_;
  wire _0637_;
  wire _0638_;
  wire _0639_;
  wire _0640_;
  wire _0641_;
  wire _0642_;
  wire _0643_;
  wire _0644_;
  wire _0645_;
  wire _0646_;
  wire [5:0] _0647_;
  wire [5:0] _0648_;
  wire [5:0] _0649_;
  wire [5:0] _0650_;
  wire [5:0] _0651_;
  wire [5:0] _0652_;
  wire [1:0] _0653_;
  wire [1:0] _0654_;
  wire [1:0] _0655_;
  wire [1:0] _0656_;
  wire [1:0] _0657_;
  wire [1:0] _0658_;
  wire _0659_;
  wire _0660_;
  wire _0661_;
  wire _0662_;
  wire [1:0] _0663_;
  wire [1:0] _0664_;
  wire _0665_;
  wire _0666_;
  wire _0667_;
  wire _0668_;
  wire _0669_;
  wire _0670_;
  wire _0671_;
  wire _0672_;
  wire _0673_;
  wire _0674_;
  wire _0675_;
  wire _0676_;
  wire _0677_;
  wire _0678_;
  wire _0679_;
  wire _0680_;
  wire _0681_;
  wire _0682_;
  wire _0683_;
  wire _0684_;
  wire _0685_;
  wire _0686_;
  wire _0687_;
  wire _0688_;
  wire _0689_;
  wire _0690_;
  wire _0691_;
  wire _0692_;
  wire _0693_;
  wire _0694_;
  wire _0695_;
  wire _0696_;
  wire _0697_;
  wire _0698_;
  wire _0699_;
  wire _0700_;
  wire _0701_;
  wire _0702_;
  wire _0703_;
  wire _0704_;
  wire _0705_;
  wire _0706_;
  wire _0707_;
  wire _0708_;
  wire _0709_;
  wire _0710_;
  wire _0711_;
  wire _0712_;
  wire _0713_;
  wire _0714_;
  wire _0715_;
  wire _0716_;
  wire _0717_;
  wire _0718_;
  wire [3:0] _0719_;
  wire [3:0] _0720_;
  wire [14:0] _0721_;
  wire _0722_;
  wire _0723_;
  wire _0724_;
  wire _0725_;
  wire _0726_;
  wire _0727_;
  wire _0728_;
  wire _0729_;
  wire _0730_;
  wire _0731_;
  wire _0732_;
  wire _0733_;
  wire _0734_;
  wire _0735_;
  wire _0736_;
  wire _0737_;
  wire _0738_;
  wire _0739_;
  wire _0740_;
  wire _0741_;
  wire _0742_;
  wire _0743_;
  wire _0744_;
  wire _0745_;
  wire _0746_;
  wire _0747_;
  wire _0748_;
  wire _0749_;
  wire _0750_;
  wire _0751_;
  wire _0752_;
  wire _0753_;
  wire _0754_;
  wire _0755_;
  wire _0756_;
  wire _0757_;
  wire _0758_;
  wire _0759_;
  wire _0760_;
  wire _0761_;
  wire _0762_;
  wire _0763_;
  wire _0764_;
  wire _0765_;
  wire _0766_;
  wire _0767_;
  wire _0768_;
  wire _0769_;
  wire _0770_;
  wire _0771_;
  wire _0772_;
  wire _0773_;
  wire _0774_;
  wire _0775_;
  wire _0776_;
  wire _0777_;
  wire _0778_;
  wire _0779_;
  wire _0780_;
  wire _0781_;
  wire _0782_;
  wire _0783_;
  wire _0784_;
  wire _0785_;
  wire _0786_;
  wire _0787_;
  wire _0788_;
  wire _0789_;
  wire _0790_;
  wire _0791_;
  wire _0792_;
  wire _0793_;
  wire _0794_;
  wire _0795_;
  wire _0796_;
  wire _0797_;
  wire _0798_;
  wire _0799_;
  wire _0800_;
  wire _0801_;
  wire _0802_;
  wire _0803_;
  wire _0804_;
  wire _0805_;
  wire _0806_;
  wire _0807_;
  wire _0808_;
  wire _0809_;
  wire _0810_;
  wire _0811_;
  wire _0812_;
  wire _0813_;
  wire _0814_;
  wire _0815_;
  wire _0816_;
  wire _0817_;
  wire _0818_;
  wire _0819_;
  wire _0820_;
  wire _0821_;
  wire _0822_;
  wire [3:0] _0823_;
  wire [3:0] _0824_;
  wire [3:0] _0825_;
  wire [3:0] _0826_;
  wire [3:0] _0827_;
  wire [3:0] _0828_;
  wire [3:0] _0829_;
  wire [3:0] _0830_;
  wire [3:0] _0831_;
  wire [2:0] _0832_;
  wire [2:0] _0833_;
  wire [2:0] _0834_;
  wire [3:0] _0835_;
  wire [3:0] _0836_;
  wire [3:0] _0837_;
  wire _0838_;
  wire _0839_;
  wire [2:0] _0840_;
  wire [2:0] _0841_;
  wire [2:0] _0842_;
  wire [3:0] _0843_;
  wire [3:0] _0844_;
  wire [3:0] _0845_;
  wire _0846_;
  wire [3:0] _0847_;
  wire [3:0] _0848_;
  wire [3:0] _0849_;
  wire _0850_;
  wire _0851_;
  wire [5:0] _0852_;
  wire [5:0] _0853_;
  wire [5:0] _0854_;
  wire [31:0] _0855_;
  wire [31:0] _0856_;
  wire [31:0] _0857_;
  wire [31:0] _0858_;
  wire [31:0] _0859_;
  wire [31:0] _0860_;
  wire [31:0] _0861_;
  wire [31:0] _0862_;
  wire [31:0] _0863_;
  wire [31:0] _0864_;
  wire [31:0] _0865_;
  wire [31:0] _0866_;
  wire [31:0] _0867_;
  wire [31:0] _0868_;
  wire [31:0] _0869_;
  wire [31:0] _0870_;
  wire [31:0] _0871_;
  wire [31:0] _0872_;
  wire [5:0] _0873_;
  wire [5:0] _0874_;
  wire [5:0] _0875_;
  wire [5:0] _0876_;
  wire [5:0] _0877_;
  wire [5:0] _0878_;
  wire [5:0] _0879_;
  wire [5:0] _0880_;
  wire [5:0] _0881_;
  wire [5:0] _0882_;
  wire [5:0] _0883_;
  wire [5:0] _0884_;
  wire [5:0] _0885_;
  wire [5:0] _0886_;
  wire [5:0] _0887_;
  wire [5:0] _0888_;
  wire [5:0] _0889_;
  wire [5:0] _0890_;
  wire [3:0] _0891_;
  wire [3:0] _0892_;
  wire [3:0] _0893_;
  wire [3:0] _0894_;
  wire [3:0] _0895_;
  wire [3:0] _0896_;
  wire [3:0] _0897_;
  wire [3:0] _0898_;
  wire [3:0] _0899_;
  wire [3:0] _0900_;
  wire [3:0] _0901_;
  wire [3:0] _0902_;
  wire _0903_;
  wire _0904_;
  wire _0905_;
  wire _0906_;
  wire _0907_;
  wire _0908_;
  wire _0909_;
  wire _0910_;
  wire _0911_;
  wire _0912_;
  wire _0913_;
  wire _0914_;
  wire _0915_;
  wire _0916_;
  wire _0917_;
  wire _0918_;
  wire _0919_;
  wire _0920_;
  wire _0921_;
  wire _0922_;
  wire [3:0] _0923_;
  wire [3:0] _0924_;
  wire [3:0] _0925_;
  wire _0926_;
  wire _0927_;
  wire [31:0] _0928_;
  wire [31:0] _0929_;
  wire [31:0] _0930_;
  wire _0931_;
  wire _0932_;
  wire _0933_;
  wire [5:0] _0934_;
  wire [5:0] _0935_;
  wire [5:0] _0936_;
  wire _0937_;
  wire _0938_;
  wire _0939_;
  wire _0940_;
  wire [1:0] _0941_;
  wire [1:0] _0942_;
  wire [1:0] _0943_;
  wire [2:0] _0944_;
  wire [2:0] _0945_;
  wire [2:0] _0946_;
  wire _0947_;
  wire _0948_;
  wire _0949_;
  wire _0950_;
  wire [2:0] _0951_;
  wire [2:0] _0952_;
  wire [2:0] _0953_;
  wire [2:0] _0954_;
  wire [2:0] _0955_;
  wire [2:0] _0956_;
  wire [5:0] _0957_;
  wire [5:0] _0958_;
  wire [5:0] _0959_;
  wire [5:0] _0960_;
  wire [5:0] _0961_;
  wire [5:0] _0962_;
  wire [5:0] _0963_;
  wire [5:0] _0964_;
  wire [5:0] _0965_;
  wire [5:0] _0966_;
  wire [5:0] _0967_;
  wire [5:0] _0968_;
  wire [5:0] _0969_;
  wire [5:0] _0970_;
  wire [5:0] _0971_;
  wire _0972_;
  wire _0973_;
  wire [3:0] _0974_;
  wire [3:0] _0975_;
  wire [3:0] _0976_;
  wire _0977_;
  wire _0978_;
  wire [3:0] _0979_;
  wire [3:0] _0980_;
  wire [3:0] _0981_;
  wire _0982_;
  wire _0983_;
  wire _0984_;
  wire [3:0] _0985_;
  wire [3:0] _0986_;
  wire [3:0] _0987_;
  wire _0988_;
  wire _0989_;
  wire _0990_;
  wire _0991_;
  wire [3:0] _0992_;
  wire [3:0] _0993_;
  wire [3:0] _0994_;
  wire [3:0] _0995_;
  wire [3:0] _0996_;
  wire [3:0] _0997_;
  wire _0998_;
  wire _0999_;
  wire [3:0] _1000_;
  wire [3:0] _1001_;
  wire [3:0] _1002_;
  wire [3:0] _1003_;
  wire [3:0] _1004_;
  wire [3:0] _1005_;
  wire [3:0] _1006_;
  wire [3:0] _1007_;
  wire [3:0] _1008_;
  wire [3:0] _1009_;
  wire [3:0] _1010_;
  wire _1011_;
  wire _1012_;
  wire [3:0] _1013_;
  wire _1014_;
  wire _1015_;
  wire _1016_;
  wire _1017_;
  wire [3:0] _1018_;
  wire [2:0] _1019_;
  wire [2:0] _1020_;
  wire [2:0] _1021_;
  wire [31:0] _1022_;
  wire [31:0] _1023_;
  wire [31:0] _1024_;
  wire _1025_;
  wire _1026_;
  wire _1027_;
  wire _1028_;
  wire _1029_;
  wire _1030_;
  wire [3:0] _1031_;
  wire [3:0] _1032_;
  wire [3:0] _1033_;
  wire [3:0] _1034_;
  wire [3:0] _1035_;
  wire [3:0] _1036_;
  wire [3:0] _1037_;
  wire [3:0] _1038_;
  wire [3:0] _1039_;
  wire [3:0] _1040_;
  wire [3:0] _1041_;
  wire [3:0] _1042_;
  wire [3:0] _1043_;
  wire [3:0] _1044_;
  wire [3:0] _1045_;
  wire [3:0] _1046_;
  wire [3:0] _1047_;
  wire [3:0] _1048_;
  wire [3:0] _1049_;
  wire [3:0] _1050_;
  wire [3:0] _1051_;
  wire [3:0] _1052_;
  wire [3:0] _1053_;
  wire [3:0] _1054_;
  wire [3:0] _1055_;
  wire [3:0] _1056_;
  wire [3:0] _1057_;
  wire [3:0] _1058_;
  wire [3:0] _1059_;
  wire [3:0] _1060_;
  wire [3:0] _1061_;
  wire [3:0] _1062_;
  wire [3:0] _1063_;
  wire [3:0] _1064_;
  wire [3:0] _1065_;
  wire [3:0] _1066_;
  wire [3:0] _1067_;
  wire [3:0] _1068_;
  wire [3:0] _1069_;
  wire [3:0] _1070_;
  wire [3:0] _1071_;
  wire [3:0] _1072_;
  wire [3:0] _1073_;
  wire [3:0] _1074_;
  wire [3:0] _1075_;
  wire [3:0] _1076_;
  wire [3:0] _1077_;
  wire _1078_;
  wire _1079_;
  wire _1080_;
  wire _1081_;
  wire _1082_;
  wire _1083_;
  wire _1084_;
  wire _1085_;
  wire [1:0] _1086_;
  wire [1:0] _1087_;
  wire [1:0] _1088_;
  wire [31:0] _1089_;
  wire [31:0] _1090_;
  wire [31:0] _1091_;
  wire [31:0] _1092_;
  wire [31:0] _1093_;
  wire [31:0] _1094_;
  wire [5:0] _1095_;
  wire [5:0] _1096_;
  wire [5:0] _1097_;
  wire _1098_;
  wire _1099_;
  wire _1100_;
  wire _1101_;
  wire _1102_;
  wire _1103_;
  wire _1104_;
  wire _1105_;
  wire _1106_;
  wire _1107_;
  wire [31:0] _1108_;
  wire _1109_;
  wire _1110_;
  wire _1111_;
  wire _1112_;
  wire _1113_;
  wire _1114_;
  wire _1115_;
  wire _1116_;
  wire _1117_;
  wire _1118_;
  wire _1119_;
  wire _1120_;
  wire _1121_;
  wire _1122_;
  wire _1123_;
  wire _1124_;
  wire _1125_;
  wire _1126_;
  wire _1127_;
  wire _1128_;
  wire _1129_;
  wire _1130_;
  wire _1131_;
  wire _1132_;
  wire _1133_;
  wire _1134_;
  wire _1135_;
  wire _1136_;
  wire [3:0] _1137_;
  wire [3:0] _1138_;
  wire [3:0] _1139_;
  wire [3:0] _1140_;
  wire [3:0] _1141_;
  wire [1:0] _1142_;
  wire [2:0] _1143_;
  wire [3:0] _1144_;
  wire [1:0] _1145_;
  wire [3:0] _1146_;
  wire [4:0] _1147_;
  wire [1:0] _1148_;
  wire _1149_;
  wire _1150_;
  wire _1151_;
  wire _1152_;
  wire _1153_;
  wire [3:0] _1154_;
  wire [3:0] _1155_;
  wire [3:0] _1156_;
  wire [3:0] _1157_;
  wire [3:0] _1158_;
  wire [3:0] _1159_;
  wire [3:0] _1160_;
  wire [3:0] _1161_;
  wire [3:0] _1162_;
  wire [3:0] _1163_;
  wire [3:0] _1164_;
  wire [3:0] _1165_;
  wire [3:0] _1166_;
  wire [3:0] _1167_;
  wire [3:0] _1168_;
  wire [3:0] _1169_;
  wire [3:0] _1170_;
  wire [3:0] _1171_;
  wire [3:0] _1172_;
  wire [3:0] _1173_;
  wire [3:0] _1174_;
  wire [3:0] _1175_;
  wire [3:0] _1176_;
  wire [3:0] _1177_;
  wire _1178_;
  wire _1179_;
  wire _1180_;
  wire _1181_;
  wire _1182_;
  wire _1183_;
  wire _1184_;
  wire _1185_;
  wire _1186_;
  wire _1187_;
  wire _1188_;
  wire [2:0] _1189_;
  wire [2:0] _1190_;
  wire [2:0] _1191_;
  wire [2:0] _1192_;
  wire [2:0] _1193_;
  wire [2:0] _1194_;
  wire [2:0] _1195_;
  wire [2:0] _1196_;
  wire [2:0] _1197_;
  wire _1198_;
  wire _1199_;
  wire _1200_;
  wire _1201_;
  wire _1202_;
  wire _1203_;
  wire _1204_;
  wire _1205_;
  wire _1206_;
  wire _1207_;
  wire _1208_;
  wire _1209_;
  wire _1210_;
  wire _1211_;
  wire _1212_;
  wire [5:0] _1213_;
  wire [5:0] _1214_;
  wire [5:0] _1215_;
  wire [5:0] _1216_;
  wire [5:0] _1217_;
  wire [5:0] _1218_;
  wire [1:0] _1219_;
  wire [1:0] _1220_;
  wire [1:0] _1221_;
  wire [1:0] _1222_;
  wire [1:0] _1223_;
  wire [1:0] _1224_;
  wire _1225_;
  wire _1226_;
  wire _1227_;
  wire _1228_;
  wire _1229_;
  wire _1230_;
  wire _1231_;
  wire _1232_;
  wire _1233_;
  wire _1234_;
  wire _1235_;
  wire _1236_;
  wire _1237_;
  wire _1238_;
  wire _1239_;
  wire _1240_;
  wire _1241_;
  wire _1242_;
  wire _1243_;
  wire _1244_;
  wire _1245_;
  wire _1246_;
  wire _1247_;
  wire _1248_;
  wire _1249_;
  wire _1250_;
  wire _1251_;
  wire _1252_;
  wire _1253_;
  wire _1254_;
  wire _1255_;
  wire _1256_;
  wire _1257_;
  wire _1258_;
  wire _1259_;
  wire _1260_;
  wire _1261_;
  wire _1262_;
  wire _1263_;
  wire _1264_;
  wire _1265_;
  wire _1266_;
  wire _1267_;
  wire _1268_;
  wire _1269_;
  wire _1270_;
  wire _1271_;
  wire _1272_;
  wire _1273_;
  wire _1274_;
  wire [3:0] _1275_;
  wire [3:0] _1276_;
  wire [3:0] _1277_;
  wire [3:0] _1278_;
  wire [3:0] _1279_;
  wire [3:0] _1280_;
  wire [3:0] _1281_;
  wire [3:0] _1282_;
  wire [3:0] _1283_;
  wire [2:0] _1284_;
  wire [2:0] _1285_;
  wire [2:0] _1286_;
  wire [3:0] _1287_;
  wire [3:0] _1288_;
  wire [3:0] _1289_;
  wire _1290_;
  wire [2:0] _1291_;
  wire [2:0] _1292_;
  wire [2:0] _1293_;
  wire [3:0] _1294_;
  wire [3:0] _1295_;
  wire [3:0] _1296_;
  wire [3:0] _1297_;
  wire [3:0] _1298_;
  wire [3:0] _1299_;
  wire _1300_;
  wire [5:0] _1301_;
  wire [5:0] _1302_;
  wire [5:0] _1303_;
  wire [31:0] _1304_;
  wire [31:0] _1305_;
  wire [31:0] _1306_;
  wire [31:0] _1307_;
  wire [31:0] _1308_;
  wire [31:0] _1309_;
  wire [31:0] _1310_;
  wire [31:0] _1311_;
  wire [31:0] _1312_;
  wire [31:0] _1313_;
  wire [31:0] _1314_;
  wire [31:0] _1315_;
  wire [31:0] _1316_;
  wire [31:0] _1317_;
  wire [31:0] _1318_;
  wire [31:0] _1319_;
  wire [31:0] _1320_;
  wire [31:0] _1321_;
  wire [5:0] _1322_;
  wire [5:0] _1323_;
  wire [5:0] _1324_;
  wire [5:0] _1325_;
  wire [5:0] _1326_;
  wire [5:0] _1327_;
  wire [5:0] _1328_;
  wire [5:0] _1329_;
  wire [5:0] _1330_;
  wire [5:0] _1331_;
  wire [5:0] _1332_;
  wire [5:0] _1333_;
  wire [5:0] _1334_;
  wire [5:0] _1335_;
  wire [5:0] _1336_;
  wire [5:0] _1337_;
  wire [5:0] _1338_;
  wire [5:0] _1339_;
  wire [3:0] _1340_;
  wire [3:0] _1341_;
  wire [3:0] _1342_;
  wire [3:0] _1343_;
  wire [3:0] _1344_;
  wire [3:0] _1345_;
  wire [3:0] _1346_;
  wire [3:0] _1347_;
  wire [3:0] _1348_;
  wire [3:0] _1349_;
  wire [3:0] _1350_;
  wire [3:0] _1351_;
  wire _1352_;
  wire _1353_;
  wire _1354_;
  wire _1355_;
  wire _1356_;
  wire _1357_;
  wire _1358_;
  wire _1359_;
  wire _1360_;
  wire _1361_;
  wire _1362_;
  wire _1363_;
  wire [3:0] _1364_;
  wire [3:0] _1365_;
  wire [3:0] _1366_;
  wire _1367_;
  wire _1368_;
  wire [31:0] _1369_;
  wire [31:0] _1370_;
  wire [31:0] _1371_;
  wire [5:0] _1372_;
  wire [5:0] _1373_;
  wire [5:0] _1374_;
  wire _1375_;
  wire [1:0] _1376_;
  wire [1:0] _1377_;
  wire [1:0] _1378_;
  wire [2:0] _1379_;
  wire [2:0] _1380_;
  wire [2:0] _1381_;
  wire [2:0] _1382_;
  wire [2:0] _1383_;
  wire [2:0] _1384_;
  wire [2:0] _1385_;
  wire [2:0] _1386_;
  wire [2:0] _1387_;
  wire [5:0] _1388_;
  wire [5:0] _1389_;
  wire [5:0] _1390_;
  wire [5:0] _1391_;
  wire [5:0] _1392_;
  wire [5:0] _1393_;
  wire [5:0] _1394_;
  wire [5:0] _1395_;
  wire [5:0] _1396_;
  wire [5:0] _1397_;
  wire [5:0] _1398_;
  wire [5:0] _1399_;
  wire _1400_;
  wire [5:0] _1401_;
  wire [5:0] _1402_;
  wire [5:0] _1403_;
  wire [3:0] _1404_;
  wire [3:0] _1405_;
  wire [3:0] _1406_;
  wire _1407_;
  wire [3:0] _1408_;
  wire [3:0] _1409_;
  wire [3:0] _1410_;
  wire _1411_;
  wire _1412_;
  wire _1413_;
  wire [3:0] _1414_;
  wire [3:0] _1415_;
  wire [3:0] _1416_;
  wire _1417_;
  wire [3:0] _1418_;
  wire [3:0] _1419_;
  wire [3:0] _1420_;
  wire [3:0] _1421_;
  wire [3:0] _1422_;
  wire [3:0] _1423_;
  wire [3:0] _1424_;
  wire [3:0] _1425_;
  wire [3:0] _1426_;
  wire [3:0] _1427_;
  wire [3:0] _1428_;
  wire [3:0] _1429_;
  wire [3:0] _1430_;
  wire [3:0] _1431_;
  wire [2:0] _1432_;
  wire [2:0] _1433_;
  wire [2:0] _1434_;
  wire [31:0] _1435_;
  wire [31:0] _1436_;
  wire [31:0] _1437_;
  wire [3:0] _1438_;
  wire [3:0] _1439_;
  wire [3:0] _1440_;
  wire [3:0] _1441_;
  wire [3:0] _1442_;
  wire [3:0] _1443_;
  wire [3:0] _1444_;
  wire [3:0] _1445_;
  wire [3:0] _1446_;
  wire [3:0] _1447_;
  wire [3:0] _1448_;
  wire [3:0] _1449_;
  wire [3:0] _1450_;
  wire [3:0] _1451_;
  wire [3:0] _1452_;
  wire [3:0] _1453_;
  wire [3:0] _1454_;
  wire [3:0] _1455_;
  wire [3:0] _1456_;
  wire [3:0] _1457_;
  wire [3:0] _1458_;
  wire [3:0] _1459_;
  wire [3:0] _1460_;
  wire [3:0] _1461_;
  wire [3:0] _1462_;
  wire [3:0] _1463_;
  wire [3:0] _1464_;
  wire [3:0] _1465_;
  wire [3:0] _1466_;
  wire [3:0] _1467_;
  wire [3:0] _1468_;
  wire [3:0] _1469_;
  wire [3:0] _1470_;
  wire [3:0] _1471_;
  wire [3:0] _1472_;
  wire [3:0] _1473_;
  wire [3:0] _1474_;
  wire [3:0] _1475_;
  wire [3:0] _1476_;
  wire [3:0] _1477_;
  wire [3:0] _1478_;
  wire [3:0] _1479_;
  wire _1480_;
  wire _1481_;
  wire _1482_;
  wire _1483_;
  wire _1484_;
  wire _1485_;
  wire _1486_;
  wire [1:0] _1487_;
  wire [1:0] _1488_;
  wire [1:0] _1489_;
  wire [31:0] _1490_;
  wire [31:0] _1491_;
  wire [31:0] _1492_;
  wire [31:0] _1493_;
  wire [31:0] _1494_;
  wire [31:0] _1495_;
  wire [5:0] _1496_;
  wire [5:0] _1497_;
  wire [5:0] _1498_;
  wire [31:0] _1499_;
  wire _1500_;
  wire _1501_;
  wire [3:0] _1502_;
  wire [3:0] _1503_;
  wire [3:0] _1504_;
  wire [3:0] _1505_;
  wire [3:0] _1506_;
  wire [3:0] _1507_;
  wire [3:0] _1508_;
  wire [3:0] _1509_;
  wire _1510_;
  wire _1511_;
  wire _1512_;
  wire _1513_;
  wire [2:0] _1514_;
  wire [2:0] _1515_;
  wire _1516_;
  wire _1517_;
  wire _1518_;
  wire _1519_;
  wire _1520_;
  wire _1521_;
  wire _1522_;
  wire [5:0] _1523_;
  wire [1:0] _1524_;
  wire _1525_;
  wire [3:0] _1526_;
  wire [3:0] _1527_;
  wire [3:0] _1528_;
  wire [2:0] _1529_;
  wire [3:0] _1530_;
  wire [31:0] _1531_;
  wire [31:0] _1532_;
  wire [31:0] _1533_;
  wire [31:0] _1534_;
  wire [31:0] _1535_;
  wire [5:0] _1536_;
  wire [5:0] _1537_;
  wire [5:0] _1538_;
  wire [5:0] _1539_;
  wire [5:0] _1540_;
  wire [3:0] _1541_;
  wire [3:0] _1542_;
  wire [3:0] _1543_;
  wire [3:0] _1544_;
  wire _1545_;
  wire _1546_;
  wire _1547_;
  wire _1548_;
  wire [3:0] _1549_;
  wire _1550_;
  wire [1:0] _1551_;
  wire [2:0] _1552_;
  wire [2:0] _1553_;
  wire [5:0] _1554_;
  wire [5:0] _1555_;
  wire [5:0] _1556_;
  wire [3:0] _1557_;
  wire [3:0] _1558_;
  wire _1559_;
  wire [3:0] _1560_;
  wire [3:0] _1561_;
  wire [3:0] _1562_;
  wire [3:0] _1563_;
  wire [3:0] _1564_;
  wire [2:0] _1565_;
  wire [3:0] _1566_;
  wire [3:0] _1567_;
  wire [3:0] _1568_;
  wire [3:0] _1569_;
  wire [3:0] _1570_;
  wire [3:0] _1571_;
  wire [3:0] _1572_;
  wire [3:0] _1573_;
  wire [3:0] _1574_;
  wire [3:0] _1575_;
  wire [3:0] _1576_;
  wire [3:0] _1577_;
  wire [3:0] _1578_;
  wire _1579_;
  wire _1580_;
  wire [31:0] _1581_;
  wire [31:0] _1582_;
  wire _1583_;
  wire _1584_;
  wire _1585_;
  wire _1586_;
  wire _1587_;
  wire _1588_;
  wire _1589_;
  wire _1590_;
  wire _1591_;
  wire _1592_;
  wire _1593_;
  wire _1594_;
  wire _1595_;
  wire _1596_;
  wire _1597_;
  wire _1598_;
  wire _1599_;
  wire _1600_;
  wire [31:0] _1601_;
  wire [31:0] _1602_;
  wire [3:0] _1603_;
  wire [3:0] _1604_;
  wire [3:0] _1605_;
  wire [3:0] _1606_;
  wire [3:0] _1607_;
  wire [3:0] _1608_;
  wire [3:0] _1609_;
  wire [3:0] _1610_;
  wire [3:0] _1611_;
  wire [3:0] _1612_;
  wire [3:0] _1613_;
  wire [3:0] _1614_;
  wire [3:0] _1615_;
  wire [3:0] _1616_;
  wire _1617_;
  wire _1618_;
  wire _1619_;
  wire _1620_;
  wire _1621_;
  wire _1622_;
  wire _1623_;
  wire _1624_;
  wire _1625_;
  wire _1626_;
  wire [2:0] _1627_;
  wire [2:0] _1628_;
  wire [2:0] _1629_;
  wire [2:0] _1630_;
  wire _1631_;
  wire _1632_;
  wire _1633_;
  wire _1634_;
  wire _1635_;
  wire _1636_;
  wire _1637_;
  wire _1638_;
  wire _1639_;
  wire _1640_;
  wire _1641_;
  wire _1642_;
  wire [5:0] _1643_;
  wire [5:0] _1644_;
  wire [1:0] _1645_;
  wire [1:0] _1646_;
  wire _1647_;
  wire _1648_;
  wire _1649_;
  wire _1650_;
  wire _1651_;
  wire _1652_;
  wire _1653_;
  wire _1654_;
  wire _1655_;
  wire _1656_;
  wire _1657_;
  wire _1658_;
  wire _1659_;
  wire _1660_;
  wire _1661_;
  wire _1662_;
  wire _1663_;
  wire _1664_;
  wire _1665_;
  wire _1666_;
  wire _1667_;
  wire _1668_;
  wire _1669_;
  wire _1670_;
  wire _1671_;
  wire _1672_;
  wire _1673_;
  wire _1674_;
  wire _1675_;
  wire _1676_;
  wire _1677_;
  wire _1678_;
  wire _1679_;
  wire _1680_;
  wire _1681_;
  wire _1682_;
  wire _1683_;
  wire _1684_;
  wire _1685_;
  wire _1686_;
  wire _1687_;
  wire _1688_;
  wire _1689_;
  wire _1690_;
  wire _1691_;
  wire _1692_;
  wire _1693_;
  wire _1694_;
  wire _1695_;
  wire _1696_;
  wire _1697_;
  wire _1698_;
  wire _1699_;
  wire _1700_;
  wire _1701_;
  wire _1702_;
  wire _1703_;
  wire _1704_;
  wire _1705_;
  wire _1706_;
  wire _1707_;
  wire _1708_;
  wire _1709_;
  wire _1710_;
  wire _1711_;
  wire _1712_;
  wire _1713_;
  wire _1714_;
  wire _1715_;
  wire _1716_;
  wire _1717_;
  wire _1718_;
  wire _1719_;
  wire [31:0] _1720_;
  wire [31:0] _1721_;
  wire [31:0] _1722_;
  wire [31:0] _1723_;
  wire [31:0] _1724_;
  wire [31:0] _1725_;
  wire [31:0] _1726_;
  wire [31:0] _1727_;
  wire [5:0] _1728_;
  wire [5:0] _1729_;
  wire [5:0] _1730_;
  wire [5:0] _1731_;
  wire [5:0] _1732_;
  wire [5:0] _1733_;
  wire [5:0] _1734_;
  wire [5:0] _1735_;
  wire [5:0] _1736_;
  wire [5:0] _1737_;
  wire [3:0] _1738_;
  wire [3:0] _1739_;
  wire [3:0] _1740_;
  wire [3:0] _1741_;
  wire [3:0] _1742_;
  wire [3:0] _1743_;
  wire _1744_;
  wire _1745_;
  wire _1746_;
  wire _1747_;
  wire _1748_;
  wire _1749_;
  wire _1750_;
  wire _1751_;
  wire _1752_;
  wire _1753_;
  wire _1754_;
  wire _1755_;
  wire _1756_;
  wire _1757_;
  wire _1758_;
  wire _1759_;
  wire _1760_;
  wire _1761_;
  wire _1762_;
  wire _1763_;
  wire _1764_;
  wire _1765_;
  wire _1766_;
  wire _1767_;
  wire _1768_;
  wire _1769_;
  wire [1:0] _1770_;
  wire [1:0] _1771_;
  wire [31:0] _1772_;
  wire [31:0] _1773_;
  wire [31:0] _1774_;
  wire [31:0] _1775_;
  wire [5:0] _1776_;
  wire [5:0] _1777_;
  input branch_not_set_i;
  wire branch_not_set_i;
  input branch_not_set_i_t0;
  wire branch_not_set_i_t0;
  input branch_set_i;
  wire branch_set_i;
  input branch_set_i_t0;
  wire branch_set_i_t0;
  input branch_set_spec_i;
  wire branch_set_spec_i;
  input branch_set_spec_i_t0;
  wire branch_set_spec_i_t0;
  input clk_i;
  wire clk_i;
  output controller_run_o;
  wire controller_run_o;
  output controller_run_o_t0;
  wire controller_run_o_t0;
  input csr_mstatus_mie_i;
  wire csr_mstatus_mie_i;
  input csr_mstatus_mie_i_t0;
  wire csr_mstatus_mie_i_t0;
  input csr_mstatus_tw_i;
  wire csr_mstatus_tw_i;
  input csr_mstatus_tw_i_t0;
  wire csr_mstatus_tw_i_t0;
  output [31:0] csr_mtval_o;
  wire [31:0] csr_mtval_o;
  output [31:0] csr_mtval_o_t0;
  wire [31:0] csr_mtval_o_t0;
  wire csr_pipe_flush;
  input csr_pipe_flush_i;
  wire csr_pipe_flush_i;
  input csr_pipe_flush_i_t0;
  wire csr_pipe_flush_i_t0;
  wire csr_pipe_flush_t0;
  output csr_restore_dret_id_o;
  wire csr_restore_dret_id_o;
  output csr_restore_dret_id_o_t0;
  wire csr_restore_dret_id_o_t0;
  output csr_restore_mret_id_o;
  wire csr_restore_mret_id_o;
  output csr_restore_mret_id_o_t0;
  wire csr_restore_mret_id_o_t0;
  output csr_save_cause_o;
  wire csr_save_cause_o;
  output csr_save_cause_o_t0;
  wire csr_save_cause_o_t0;
  output csr_save_id_o;
  wire csr_save_id_o;
  output csr_save_id_o_t0;
  wire csr_save_id_o_t0;
  output csr_save_if_o;
  wire csr_save_if_o;
  output csr_save_if_o_t0;
  wire csr_save_if_o_t0;
  output csr_save_wb_o;
  wire csr_save_wb_o;
  output csr_save_wb_o_t0;
  wire csr_save_wb_o_t0;
  output ctrl_busy_o;
  wire ctrl_busy_o;
  output ctrl_busy_o_t0;
  wire ctrl_busy_o_t0;
  reg [3:0] ctrl_fsm_cs;
  reg [3:0] ctrl_fsm_cs_t0;
  wire [3:0] ctrl_fsm_ns;
  wire [3:0] ctrl_fsm_ns_t0;
  output [2:0] debug_cause_o;
  wire [2:0] debug_cause_o;
  output [2:0] debug_cause_o_t0;
  wire [2:0] debug_cause_o_t0;
  output debug_csr_save_o;
  wire debug_csr_save_o;
  output debug_csr_save_o_t0;
  wire debug_csr_save_o_t0;
  input debug_ebreakm_i;
  wire debug_ebreakm_i;
  input debug_ebreakm_i_t0;
  wire debug_ebreakm_i_t0;
  input debug_ebreaku_i;
  wire debug_ebreaku_i;
  input debug_ebreaku_i_t0;
  wire debug_ebreaku_i_t0;
  wire debug_mode_d;
  wire debug_mode_d_t0;
  output debug_mode_o;
  reg debug_mode_o;
  output debug_mode_o_t0;
  reg debug_mode_o_t0;
  input debug_req_i;
  wire debug_req_i;
  input debug_req_i_t0;
  wire debug_req_i_t0;
  input debug_single_step_i;
  wire debug_single_step_i;
  input debug_single_step_i_t0;
  wire debug_single_step_i_t0;
  wire do_single_step_d;
  wire do_single_step_d_t0;
  reg do_single_step_q;
  reg do_single_step_q_t0;
  wire dret_insn;
  input dret_insn_i;
  wire dret_insn_i;
  input dret_insn_i_t0;
  wire dret_insn_i_t0;
  wire dret_insn_t0;
  wire ebreak_into_debug;
  wire ebreak_into_debug_t0;
  wire ebrk_insn;
  input ebrk_insn_i;
  wire ebrk_insn_i;
  input ebrk_insn_i_t0;
  wire ebrk_insn_i_t0;
  wire ebrk_insn_prio;
  wire ebrk_insn_prio_t0;
  wire ebrk_insn_t0;
  wire ecall_insn;
  input ecall_insn_i;
  wire ecall_insn_i;
  input ecall_insn_i_t0;
  wire ecall_insn_i_t0;
  wire ecall_insn_prio;
  wire ecall_insn_prio_t0;
  wire ecall_insn_t0;
  wire enter_debug_mode;
  wire enter_debug_mode_prio_d;
  wire enter_debug_mode_prio_d_t0;
  reg enter_debug_mode_prio_q;
  reg enter_debug_mode_prio_q_t0;
  wire enter_debug_mode_t0;
  output [5:0] exc_cause_o;
  wire [5:0] exc_cause_o;
  output [5:0] exc_cause_o_t0;
  wire [5:0] exc_cause_o_t0;
  output [1:0] exc_pc_mux_o;
  wire [1:0] exc_pc_mux_o;
  output [1:0] exc_pc_mux_o_t0;
  wire [1:0] exc_pc_mux_o_t0;
  wire exc_req_d;
  wire exc_req_d_t0;
  wire exc_req_lsu;
  wire exc_req_lsu_t0;
  reg exc_req_q;
  reg exc_req_q_t0;
  output flush_id_o;
  wire flush_id_o;
  output flush_id_o_t0;
  wire flush_id_o_t0;
  wire halt_if;
  wire halt_if_t0;
  wire handle_irq;
  wire handle_irq_t0;
  output id_in_ready_o;
  wire id_in_ready_o;
  output id_in_ready_o_t0;
  wire id_in_ready_o_t0;
  wire id_wb_pending;
  wire id_wb_pending_t0;
  wire illegal_dret;
  wire illegal_dret_t0;
  wire illegal_insn_d;
  wire illegal_insn_d_t0;
  input illegal_insn_i;
  wire illegal_insn_i;
  input illegal_insn_i_t0;
  wire illegal_insn_i_t0;
  wire illegal_insn_prio;
  wire illegal_insn_prio_t0;
  reg illegal_insn_q;
  reg illegal_insn_q_t0;
  wire illegal_umode;
  wire illegal_umode_t0;
  input instr_bp_taken_i;
  wire instr_bp_taken_i;
  input instr_bp_taken_i_t0;
  wire instr_bp_taken_i_t0;
  input [15:0] instr_compressed_i;
  wire [15:0] instr_compressed_i;
  input [15:0] instr_compressed_i_t0;
  wire [15:0] instr_compressed_i_t0;
  wire instr_fetch_err;
  input instr_fetch_err_i;
  wire instr_fetch_err_i;
  input instr_fetch_err_i_t0;
  wire instr_fetch_err_i_t0;
  input instr_fetch_err_plus2_i;
  wire instr_fetch_err_plus2_i;
  input instr_fetch_err_plus2_i_t0;
  wire instr_fetch_err_plus2_i_t0;
  wire instr_fetch_err_prio;
  wire instr_fetch_err_prio_t0;
  wire instr_fetch_err_t0;
  input [31:0] instr_i;
  wire [31:0] instr_i;
  input [31:0] instr_i_t0;
  wire [31:0] instr_i_t0;
  input instr_is_compressed_i;
  wire instr_is_compressed_i;
  input instr_is_compressed_i_t0;
  wire instr_is_compressed_i_t0;
  output instr_req_o;
  wire instr_req_o;
  output instr_req_o_t0;
  wire instr_req_o_t0;
  output instr_valid_clear_o;
  wire instr_valid_clear_o;
  output instr_valid_clear_o_t0;
  wire instr_valid_clear_o_t0;
  input instr_valid_i;
  wire instr_valid_i;
  input instr_valid_i_t0;
  wire instr_valid_i_t0;
  input irq_nm_i;
  wire irq_nm_i;
  input irq_nm_i_t0;
  wire irq_nm_i_t0;
  input irq_pending_i;
  wire irq_pending_i;
  input irq_pending_i_t0;
  wire irq_pending_i_t0;
  input [17:0] irqs_i;
  wire [17:0] irqs_i;
  input [17:0] irqs_i_t0;
  wire [17:0] irqs_i_t0;
  input jump_set_i;
  wire jump_set_i;
  input jump_set_i_t0;
  wire jump_set_i_t0;
  input load_err_i;
  wire load_err_i;
  input load_err_i_t0;
  wire load_err_i_t0;
  wire load_err_prio;
  wire load_err_prio_t0;
  reg load_err_q;
  reg load_err_q_t0;
  input [31:0] lsu_addr_last_i;
  wire [31:0] lsu_addr_last_i;
  input [31:0] lsu_addr_last_i_t0;
  wire [31:0] lsu_addr_last_i_t0;
  wire [3:0] mfip_id;
  wire [3:0] mfip_id_t0;
  wire mret_insn;
  input mret_insn_i;
  wire mret_insn_i;
  input mret_insn_i_t0;
  wire mret_insn_i_t0;
  wire mret_insn_t0;
  wire nmi_mode_d;
  wire nmi_mode_d_t0;
  output nmi_mode_o;
  reg nmi_mode_o;
  output nmi_mode_o_t0;
  reg nmi_mode_o_t0;
  output nt_branch_mispredict_o;
  wire nt_branch_mispredict_o;
  output nt_branch_mispredict_o_t0;
  wire nt_branch_mispredict_o_t0;
  input [31:0] pc_id_i;
  wire [31:0] pc_id_i;
  input [31:0] pc_id_i_t0;
  wire [31:0] pc_id_i_t0;
  output [2:0] pc_mux_o;
  wire [2:0] pc_mux_o;
  output [2:0] pc_mux_o_t0;
  wire [2:0] pc_mux_o_t0;
  output pc_set_o;
  wire pc_set_o;
  output pc_set_o_t0;
  wire pc_set_o_t0;
  output pc_set_spec_o;
  wire pc_set_spec_o;
  output pc_set_spec_o_t0;
  wire pc_set_spec_o_t0;
  output perf_jump_o;
  wire perf_jump_o;
  output perf_jump_o_t0;
  wire perf_jump_o_t0;
  output perf_tbranch_o;
  wire perf_tbranch_o;
  output perf_tbranch_o_t0;
  wire perf_tbranch_o_t0;
  input [1:0] priv_mode_i;
  wire [1:0] priv_mode_i;
  input [1:0] priv_mode_i_t0;
  wire [1:0] priv_mode_i_t0;
  input ready_wb_i;
  wire ready_wb_i;
  input ready_wb_i_t0;
  wire ready_wb_i_t0;
  wire retain_id;
  wire retain_id_t0;
  input rst_ni;
  wire rst_ni;
  wire special_req;
  wire special_req_flush_only;
  wire special_req_flush_only_t0;
  wire special_req_pc_change;
  wire special_req_pc_change_t0;
  wire special_req_t0;
  wire stall;
  input stall_id_i;
  wire stall_id_i;
  input stall_id_i_t0;
  wire stall_id_i_t0;
  wire stall_t0;
  input stall_wb_i;
  wire stall_wb_i;
  input stall_wb_i_t0;
  wire stall_wb_i_t0;
  input store_err_i;
  wire store_err_i;
  input store_err_i_t0;
  wire store_err_i_t0;
  wire store_err_prio;
  reg store_err_prio_t0;
  reg store_err_q;
  input trigger_match_i;
  wire trigger_match_i;
  input trigger_match_i_t0;
  wire trigger_match_i_t0;
  output wb_exception_o;
  wire wb_exception_o;
  output wb_exception_o_t0;
  wire wb_exception_o_t0;
  wire wfi_insn;
  input wfi_insn_i;
  wire wfi_insn_i;
  input wfi_insn_i_t0;
  wire wfi_insn_i_t0;
  wire wfi_insn_t0;
  assign _0179_ = pc_id_i + 32'd2;
  assign ecall_insn = ecall_insn_i & instr_valid_i;
  assign mret_insn = mret_insn_i & instr_valid_i;
  assign dret_insn = dret_insn_i & instr_valid_i;
  assign wfi_insn = wfi_insn_i & instr_valid_i;
  assign ebrk_insn = ebrk_insn_i & instr_valid_i;
  assign csr_pipe_flush = csr_pipe_flush_i & instr_valid_i;
  assign instr_fetch_err = instr_fetch_err_i & instr_valid_i;
  assign illegal_dret = dret_insn & _0284_;
  assign _0181_ = csr_mstatus_tw_i & wfi_insn;
  assign illegal_umode = _1687_ & _1695_;
  assign illegal_insn_d = _1699_ & _1688_;
  assign exc_req_d = _1705_ & _1688_;
  assign _0183_ = _0284_ & debug_single_step_i;
  assign enter_debug_mode_prio_d = _1713_ & _0284_;
  assign _0185_ = trigger_match_i & _0284_;
  assign _0187_ = _0284_ & _1691_;
  assign _0189_ = irq_pending_i & csr_mstatus_mie_i;
  assign handle_irq = _0187_ & _1715_;
  assign _0191_ = _0292_ & _1692_;
  assign id_in_ready_o = _0191_ & _0334_;
  assign _0230_ = ~ pc_id_i_t0;
  assign _0462_ = pc_id_i & _0230_;
  assign _1601_ = _0462_ + 32'd2;
  assign _1108_ = pc_id_i | pc_id_i_t0;
  assign _1602_ = _1108_ + 32'd2;
  assign _1499_ = _1601_ ^ _1602_;
  assign _0180_ = _1499_ | pc_id_i_t0;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) load_err_q_t0 <= 1'h0;
    else load_err_q_t0 <= load_err_i_t0;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) store_err_prio_t0 <= 1'h0;
    else store_err_prio_t0 <= store_err_i_t0;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) exc_req_q_t0 <= 1'h0;
    else exc_req_q_t0 <= exc_req_d_t0;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) illegal_insn_q_t0 <= 1'h0;
    else illegal_insn_q_t0 <= illegal_insn_d_t0;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) do_single_step_q_t0 <= 1'h0;
    else do_single_step_q_t0 <= do_single_step_d_t0;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) enter_debug_mode_prio_q_t0 <= 1'h0;
    else enter_debug_mode_prio_q_t0 <= enter_debug_mode_prio_d_t0;
  assign _0231_ = ~ _0213_;
  assign _0232_ = ~ _0215_;
  assign _0233_ = ~ _0217_;
  assign _1500_ = debug_mode_d ^ debug_mode_o;
  assign _1501_ = nmi_mode_d ^ nmi_mode_o;
  assign _1502_ = ctrl_fsm_ns ^ ctrl_fsm_cs;
  assign _1129_ = debug_mode_d_t0 | debug_mode_o_t0;
  assign _1133_ = nmi_mode_d_t0 | nmi_mode_o_t0;
  assign _1137_ = ctrl_fsm_ns_t0 | ctrl_fsm_cs_t0;
  assign _1130_ = _1500_ | _1129_;
  assign _1134_ = _1501_ | _1133_;
  assign _1138_ = _1502_ | _1137_;
  assign _0523_ = _0213_ & debug_mode_d_t0;
  assign _0526_ = _0215_ & nmi_mode_d_t0;
  assign _0529_ = { _0217_, _0217_, _0217_, _0217_ } & ctrl_fsm_ns_t0;
  assign _0524_ = _0231_ & debug_mode_o_t0;
  assign _0527_ = _0232_ & nmi_mode_o_t0;
  assign _0530_ = { _0233_, _0233_, _0233_, _0233_ } & ctrl_fsm_cs_t0;
  assign _0525_ = _1130_ & _0214_;
  assign _0528_ = _1134_ & _0216_;
  assign _0531_ = _1138_ & { _0218_, _0218_, _0218_, _0218_ };
  assign _1131_ = _0523_ | _0524_;
  assign _1135_ = _0526_ | _0527_;
  assign _1139_ = _0529_ | _0530_;
  assign _1132_ = _1131_ | _0525_;
  assign _1136_ = _1135_ | _0528_;
  assign _1140_ = _1139_ | _0531_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) debug_mode_o_t0 <= 1'h0;
    else debug_mode_o_t0 <= _1132_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) nmi_mode_o_t0 <= 1'h0;
    else nmi_mode_o_t0 <= _1136_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) ctrl_fsm_cs_t0 <= 4'h0;
    else ctrl_fsm_cs_t0 <= _1140_;
  assign _0463_ = ecall_insn_i_t0 & instr_valid_i;
  assign _0466_ = mret_insn_i_t0 & instr_valid_i;
  assign _0469_ = dret_insn_i_t0 & instr_valid_i;
  assign _0472_ = wfi_insn_i_t0 & instr_valid_i;
  assign _0475_ = ebrk_insn_i_t0 & instr_valid_i;
  assign _0478_ = csr_pipe_flush_i_t0 & instr_valid_i;
  assign _0481_ = instr_fetch_err_i_t0 & instr_valid_i;
  assign _0484_ = dret_insn_t0 & _0284_;
  assign _0487_ = csr_mstatus_tw_i_t0 & wfi_insn;
  assign _0490_ = _1649_ & _1695_;
  assign _0493_ = _1700_ & _1688_;
  assign _0496_ = _1706_ & _1688_;
  assign _0499_ = debug_mode_o_t0 & debug_single_step_i;
  assign _0502_ = _1714_ & _0284_;
  assign _0505_ = trigger_match_i_t0 & _0284_;
  assign _0508_ = debug_mode_o_t0 & _1691_;
  assign _0511_ = irq_pending_i_t0 & csr_mstatus_mie_i;
  assign _0514_ = _0188_ & _1715_;
  assign _0517_ = stall_t0 & _1692_;
  assign _0520_ = _0192_ & _0334_;
  assign _0464_ = instr_valid_i_t0 & ecall_insn_i;
  assign _0467_ = instr_valid_i_t0 & mret_insn_i;
  assign _0470_ = instr_valid_i_t0 & dret_insn_i;
  assign _0473_ = instr_valid_i_t0 & wfi_insn_i;
  assign _0476_ = instr_valid_i_t0 & ebrk_insn_i;
  assign _0479_ = instr_valid_i_t0 & csr_pipe_flush_i;
  assign _0482_ = instr_valid_i_t0 & instr_fetch_err_i;
  assign _0485_ = debug_mode_o_t0 & dret_insn;
  assign _0488_ = wfi_insn_t0 & csr_mstatus_tw_i;
  assign _0491_ = _1696_ & _1687_;
  assign _0494_ = _1141_[3] & _1699_;
  assign _0497_ = _1141_[3] & _1705_;
  assign _0500_ = debug_single_step_i_t0 & _0284_;
  assign _0503_ = debug_mode_o_t0 & _1713_;
  assign _0506_ = debug_mode_o_t0 & trigger_match_i;
  assign _0509_ = nmi_mode_o_t0 & _0284_;
  assign _0512_ = csr_mstatus_mie_i_t0 & irq_pending_i;
  assign _0515_ = _1716_ & _0187_;
  assign _0518_ = halt_if_t0 & _0292_;
  assign _0521_ = retain_id_t0 & _0191_;
  assign _0465_ = ecall_insn_i_t0 & instr_valid_i_t0;
  assign _0468_ = mret_insn_i_t0 & instr_valid_i_t0;
  assign _0471_ = dret_insn_i_t0 & instr_valid_i_t0;
  assign _0474_ = wfi_insn_i_t0 & instr_valid_i_t0;
  assign _0477_ = ebrk_insn_i_t0 & instr_valid_i_t0;
  assign _0480_ = csr_pipe_flush_i_t0 & instr_valid_i_t0;
  assign _0483_ = instr_fetch_err_i_t0 & instr_valid_i_t0;
  assign _0486_ = dret_insn_t0 & debug_mode_o_t0;
  assign _0489_ = csr_mstatus_tw_i_t0 & wfi_insn_t0;
  assign _0492_ = _1649_ & _1696_;
  assign _0495_ = _1700_ & _1141_[3];
  assign _0498_ = _1706_ & _1141_[3];
  assign _0501_ = debug_mode_o_t0 & debug_single_step_i_t0;
  assign _0504_ = _1714_ & debug_mode_o_t0;
  assign _0507_ = trigger_match_i_t0 & debug_mode_o_t0;
  assign _0510_ = debug_mode_o_t0 & nmi_mode_o_t0;
  assign _0513_ = irq_pending_i_t0 & csr_mstatus_mie_i_t0;
  assign _0516_ = _0188_ & _1716_;
  assign _0519_ = stall_t0 & halt_if_t0;
  assign _0522_ = _0192_ & retain_id_t0;
  assign _1109_ = _0463_ | _0464_;
  assign _1110_ = _0466_ | _0467_;
  assign _1111_ = _0469_ | _0470_;
  assign _1112_ = _0472_ | _0473_;
  assign _1113_ = _0475_ | _0476_;
  assign _1114_ = _0478_ | _0479_;
  assign _1115_ = _0481_ | _0482_;
  assign _1116_ = _0484_ | _0485_;
  assign _1117_ = _0487_ | _0488_;
  assign _1118_ = _0490_ | _0491_;
  assign _1119_ = _0493_ | _0494_;
  assign _1120_ = _0496_ | _0497_;
  assign _1121_ = _0499_ | _0500_;
  assign _1122_ = _0502_ | _0503_;
  assign _1123_ = _0505_ | _0506_;
  assign _1124_ = _0508_ | _0509_;
  assign _1125_ = _0511_ | _0512_;
  assign _1126_ = _0514_ | _0515_;
  assign _1127_ = _0517_ | _0518_;
  assign _1128_ = _0520_ | _0521_;
  assign ecall_insn_t0 = _1109_ | _0465_;
  assign mret_insn_t0 = _1110_ | _0468_;
  assign dret_insn_t0 = _1111_ | _0471_;
  assign wfi_insn_t0 = _1112_ | _0474_;
  assign ebrk_insn_t0 = _1113_ | _0477_;
  assign csr_pipe_flush_t0 = _1114_ | _0480_;
  assign instr_fetch_err_t0 = _1115_ | _0483_;
  assign illegal_dret_t0 = _1116_ | _0486_;
  assign _0182_ = _1117_ | _0489_;
  assign illegal_umode_t0 = _1118_ | _0492_;
  assign illegal_insn_d_t0 = _1119_ | _0495_;
  assign exc_req_d_t0 = _1120_ | _0498_;
  assign _0184_ = _1121_ | _0501_;
  assign enter_debug_mode_prio_d_t0 = _1122_ | _0504_;
  assign _0186_ = _1123_ | _0507_;
  assign _0188_ = _1124_ | _0510_;
  assign _0190_ = _1125_ | _0513_;
  assign handle_irq_t0 = _1126_ | _0516_;
  assign _0192_ = _1127_ | _0519_;
  assign id_in_ready_o_t0 = _1128_ | _0522_;
  assign _0428_ = | { _1141_[3:2], dret_insn_t0, mret_insn_t0 };
  assign _0430_ = | _1141_[3:2];
  assign _0429_ = | { _1141_[3:2], mret_insn_t0 };
  assign _0432_ = | { _1142_[1], handle_irq_t0 };
  assign _0433_ = | { _1143_[1], _1142_[1], handle_irq_t0 };
  assign _0435_ = | { _1144_[3], enter_debug_mode_t0, handle_irq_t0, id_in_ready_o_t0 };
  assign _0436_ = | { _0040_, _1145_[1] };
  assign _0447_ = | priv_mode_i_t0;
  assign _0234_ = ~ { _1141_[3:2], dret_insn_t0, mret_insn_t0 };
  assign _0236_ = ~ _1141_[3:2];
  assign _0235_ = ~ { _1141_[3:2], mret_insn_t0 };
  assign _0238_ = ~ { _1142_[1], handle_irq_t0 };
  assign _0239_ = ~ { _1142_[1], _1143_[1], handle_irq_t0 };
  assign _0241_ = ~ { _1144_[3], id_in_ready_o_t0, handle_irq_t0, enter_debug_mode_t0 };
  assign _0242_ = ~ { _1145_[1], _0040_ };
  assign _0278_ = ~ priv_mode_i_t0;
  assign _0298_ = ~ ctrl_fsm_cs_t0;
  assign _0532_ = { _1719_, _1686_, dret_insn, mret_insn } & _0234_;
  assign _0536_ = { _1719_, _1686_ } & _0236_;
  assign _0534_ = { _1719_, _1686_, mret_insn } & _0235_;
  assign _0540_ = { _1759_, handle_irq } & _0238_;
  assign _0542_ = { _1759_, _1657_, handle_irq } & _0239_;
  assign _0545_ = { _1761_, id_in_ready_o, handle_irq, enter_debug_mode } & _0241_;
  assign _0547_ = { _1762_, _1677_ } & _0242_;
  assign _0663_ = priv_mode_i & _0278_;
  assign _0719_ = ctrl_fsm_cs & _0298_;
  assign _0533_ = 4'h8 & _0234_;
  assign _0535_ = 3'h5 & _0235_;
  assign _0537_ = 2'h3 & _0236_;
  assign _0539_ = 3'h4 & _0235_;
  assign _0541_ = 2'h2 & _0238_;
  assign _0543_ = 3'h5 & _0239_;
  assign _0546_ = 4'h8 & _0241_;
  assign _0548_ = 2'h2 & _0242_;
  assign _0664_ = 2'h3 & _0278_;
  assign _1010_ = 4'h1 & _0298_;
  assign _1013_ = 4'h4 & _0298_;
  assign _1018_ = 4'h5 & _0298_;
  assign _1031_ = 4'h7 & _0298_;
  assign _0720_ = 4'h6 & _0298_;
  assign _1032_ = 4'h9 & _0298_;
  assign _1033_ = 4'h8 & _0298_;
  assign _1034_ = 4'h3 & _0298_;
  assign _1035_ = 4'h2 & _0298_;
  assign _1583_ = _0532_ == _0533_;
  assign _1584_ = _0534_ == _0535_;
  assign _1585_ = _0536_ == _0537_;
  assign _1586_ = _0534_ == _0539_;
  assign _1587_ = _0540_ == _0541_;
  assign _1588_ = _0542_ == _0543_;
  assign _1589_ = _0545_ == _0546_;
  assign _1590_ = _0547_ == _0548_;
  assign _1591_ = _0663_ == _0664_;
  assign _1593_ = _0719_ == _1010_;
  assign _1594_ = _0719_ == _1013_;
  assign _1595_ = _0719_ == _1018_;
  assign _1596_ = _0719_ == _1031_;
  assign _1592_ = _0719_ == _0720_;
  assign _1597_ = _0719_ == _1032_;
  assign _1598_ = _0719_ == _1033_;
  assign _1599_ = _0719_ == _1034_;
  assign _1600_ = _0719_ == _1035_;
  assign _0194_ = _1583_ & _0428_;
  assign _0196_ = _1584_ & _0429_;
  assign _0198_ = _1585_ & _0430_;
  assign _0202_ = _1586_ & _0429_;
  assign _0204_ = _1587_ & _0432_;
  assign _0206_ = _1588_ & _0433_;
  assign _0210_ = _1589_ & _0435_;
  assign _0212_ = _1590_ & _0436_;
  assign _1649_ = _1591_ & _0447_;
  assign _1765_ = _1593_ & _0448_;
  assign _1144_[3] = _1594_ & _0448_;
  assign controller_run_o_t0 = _1595_ & _0448_;
  assign _1142_[1] = _1596_ & _0448_;
  assign _1141_[3] = _1592_ & _0448_;
  assign _1757_ = _1597_ & _0448_;
  assign _0630_ = _1598_ & _0448_;
  assign _1145_[1] = _1599_ & _0448_;
  assign _0659_ = _1600_ & _0448_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) debug_mode_o <= 1'h0;
    else if (_0213_) debug_mode_o <= debug_mode_d;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) nmi_mode_o <= 1'h0;
    else if (_0215_) nmi_mode_o <= nmi_mode_d;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) ctrl_fsm_cs <= 4'h0;
    else if (_0217_) ctrl_fsm_cs <= ctrl_fsm_ns;
  assign _0665_ = _1681_ & _1682_;
  assign _0668_ = stall_t0 & _1666_;
  assign _0671_ = _1654_ & _1667_;
  assign _0674_ = irq_nm_i_t0 & _1668_;
  assign _0677_ = ebreak_into_debug_t0 & _1669_;
  assign _0680_ = csr_pipe_flush_t0 & handle_irq;
  assign _0683_ = ebrk_insn_prio_t0 & ebreak_into_debug;
  assign _0686_ = enter_debug_mode_prio_q_t0 & _1670_;
  assign _0666_ = _1683_ & _1680_;
  assign _0669_ = special_req_t0 & _1665_;
  assign _0672_ = id_wb_pending_t0 & _1653_;
  assign _0675_ = nmi_mode_o_t0 & irq_nm_i;
  assign _0678_ = debug_mode_o_t0 & ebreak_into_debug;
  assign _0681_ = handle_irq_t0 & csr_pipe_flush;
  assign _0684_ = ebreak_into_debug_t0 & ebrk_insn_prio;
  assign _0687_ = _1662_ & enter_debug_mode_prio_q;
  assign _0667_ = _1681_ & _1683_;
  assign _0670_ = stall_t0 & special_req_t0;
  assign _0673_ = _1654_ & id_wb_pending_t0;
  assign _0676_ = irq_nm_i_t0 & nmi_mode_o_t0;
  assign _0682_ = csr_pipe_flush_t0 & handle_irq_t0;
  assign _0685_ = ebrk_insn_prio_t0 & ebreak_into_debug_t0;
  assign _0688_ = enter_debug_mode_prio_q_t0 & _1662_;
  assign _1228_ = _0665_ | _0666_;
  assign _1229_ = _0668_ | _0669_;
  assign _1230_ = _0671_ | _0672_;
  assign _1231_ = _0674_ | _0675_;
  assign _1232_ = _0677_ | _0678_;
  assign _1233_ = _0680_ | _0681_;
  assign _1234_ = _0683_ | _0684_;
  assign _1235_ = _0686_ | _0687_;
  assign _0123_ = _1228_ | _0667_;
  assign _1654_ = _1229_ | _0670_;
  assign _1656_ = _1230_ | _0673_;
  assign _1143_[1] = _1231_ | _0676_;
  assign _0036_ = _1232_ | _0679_;
  assign _1660_ = _1233_ | _0682_;
  assign _1662_ = _1234_ | _0685_;
  assign _1664_ = _1235_ | _0688_;
  assign _0431_ = | { _0220_, _1141_[3] };
  assign _0434_ = | { _1142_[1], _1141_[3] };
  assign _0440_ = | { _0630_, _1767_, _1765_, _1757_ };
  assign _0441_ = | { _0659_, _0630_, _1757_, _1145_[1] };
  assign _0442_ = | { _0630_, _1765_, _1757_, _1144_[3], _1142_[1], _1141_[3], controller_run_o_t0 };
  assign _0443_ = | { _0630_, _1757_, _1142_[1] };
  assign _0444_ = | { _0659_, _1145_[1], _1141_[3] };
  assign _0445_ = | { _0630_, _1757_ };
  assign _0446_ = | { _1099_, _1144_[3], controller_run_o_t0 };
  assign _0449_ = | irqs_i_t0[14:0];
  assign _0448_ = | ctrl_fsm_cs_t0;
  assign _0237_ = ~ { _0220_, _1141_[3] };
  assign _0240_ = ~ { _1141_[3], _1142_[1] };
  assign _0243_ = ~ { _1767_, _1765_, _0630_, _1757_ };
  assign _0244_ = ~ { _0659_, _1145_[1], _0630_, _1757_ };
  assign _0245_ = ~ { _1765_, _1144_[3], controller_run_o_t0, _1142_[1], _0630_, _1757_, _1141_[3] };
  assign _0246_ = ~ { _1142_[1], _0630_, _1757_ };
  assign _0247_ = ~ { _0659_, _1145_[1], _1141_[3] };
  assign _0248_ = ~ { _0630_, _1757_ };
  assign _0257_ = ~ { _1144_[3], controller_run_o_t0, _1099_ };
  assign _0299_ = ~ irqs_i_t0[14:0];
  assign _0538_ = { _0219_, _1719_ } & _0237_;
  assign _0544_ = { _1719_, _1759_ } & _0240_;
  assign _0549_ = { _1766_, _1764_, _1758_, _1756_ } & _0243_;
  assign _0550_ = { _1763_, _1762_, _1758_, _1756_ } & _0244_;
  assign _0551_ = { _1764_, _1761_, _1760_, _1759_, _1758_, _1756_, _1719_ } & _0245_;
  assign _0552_ = { _1759_, _1758_, _1756_ } & _0246_;
  assign _0553_ = { _1763_, _1762_, _1719_ } & _0247_;
  assign _0554_ = { _1758_, _1756_ } & _0248_;
  assign _0570_ = { _1761_, _1760_, _1098_ } & _0257_;
  assign _0721_ = irqs_i[14:0] & _0299_;
  assign _0450_ = ! _0538_;
  assign _0451_ = ! _0544_;
  assign _0452_ = ! _0549_;
  assign _0453_ = ! _0550_;
  assign _0454_ = ! _0551_;
  assign _0455_ = ! _0552_;
  assign _0456_ = ! _0553_;
  assign _0457_ = ! _0554_;
  assign _0458_ = ! _0570_;
  assign _0459_ = ! _0663_;
  assign _0460_ = ! _0721_;
  assign _0461_ = ! _0719_;
  assign _0200_ = _0450_ & _0431_;
  assign _0208_ = _0451_ & _0434_;
  assign _0222_ = _0452_ & _0440_;
  assign _0224_ = _0453_ & _0441_;
  assign instr_req_o_t0 = _0454_ & _0442_;
  assign _0226_ = _0455_ & _0443_;
  assign _0229_ = _0456_ & _0444_;
  assign _0220_ = _0457_ & _0445_;
  assign _0427_ = _0458_ & _0446_;
  assign _1651_ = _0459_ & _0447_;
  assign _1690_ = _0460_ & _0449_;
  assign _1767_ = _0461_ & _0448_;
  assign _0281_ = ~ _1671_;
  assign _0283_ = ~ _1673_;
  assign _0285_ = ~ _1675_;
  assign _0287_ = ~ branch_set_i;
  assign _0289_ = ~ branch_set_spec_i;
  assign _0294_ = ~ exc_req_q;
  assign _0296_ = ~ _1684_;
  assign _0280_ = ~ irq_pending_i;
  assign _0286_ = ~ debug_single_step_i;
  assign _0288_ = ~ jump_set_i;
  assign _0293_ = ~ id_wb_pending;
  assign _0689_ = irq_nm_i_t0 & _0280_;
  assign _0692_ = _1672_ & _0282_;
  assign _0695_ = _1674_ & _0284_;
  assign _0698_ = _1676_ & _0286_;
  assign _0701_ = branch_set_i_t0 & _0288_;
  assign _0704_ = branch_set_spec_i_t0 & _0288_;
  assign _0707_ = enter_debug_mode_t0 & _0291_;
  assign _0710_ = stall_t0 & _0293_;
  assign _0713_ = exc_req_q_t0 & _0295_;
  assign _0716_ = _1685_ & _0297_;
  assign _0690_ = irq_pending_i_t0 & _0279_;
  assign _0693_ = debug_req_i_t0 & _0281_;
  assign _0696_ = debug_mode_o_t0 & _0283_;
  assign _0699_ = debug_single_step_i_t0 & _0285_;
  assign _0702_ = jump_set_i_t0 & _0287_;
  assign _0705_ = jump_set_i_t0 & _0289_;
  assign _0708_ = handle_irq_t0 & _0290_;
  assign _0711_ = id_wb_pending_t0 & _0292_;
  assign _0714_ = store_err_prio_t0 & _0294_;
  assign _0717_ = load_err_q_t0 & _0296_;
  assign _0691_ = irq_nm_i_t0 & irq_pending_i_t0;
  assign _0694_ = _1672_ & debug_req_i_t0;
  assign _0697_ = _1674_ & debug_mode_o_t0;
  assign _0700_ = _1676_ & debug_single_step_i_t0;
  assign _0703_ = branch_set_i_t0 & jump_set_i_t0;
  assign _0706_ = branch_set_spec_i_t0 & jump_set_i_t0;
  assign _0709_ = enter_debug_mode_t0 & handle_irq_t0;
  assign _0712_ = stall_t0 & id_wb_pending_t0;
  assign _0715_ = exc_req_q_t0 & store_err_prio_t0;
  assign _0718_ = _1685_ & load_err_q_t0;
  assign _1236_ = _0689_ | _0690_;
  assign _1237_ = _0692_ | _0693_;
  assign _1238_ = _0695_ | _0696_;
  assign _1239_ = _0698_ | _0699_;
  assign _1240_ = _0701_ | _0702_;
  assign _1241_ = _0704_ | _0705_;
  assign _1242_ = _0707_ | _0708_;
  assign _1243_ = _0710_ | _0711_;
  assign _1244_ = _0713_ | _0714_;
  assign _1245_ = _0716_ | _0717_;
  assign _1672_ = _1236_ | _0691_;
  assign _1674_ = _1237_ | _0694_;
  assign _1676_ = _1238_ | _0697_;
  assign _0040_ = _1239_ | _0700_;
  assign _0067_ = _1240_ | _0703_;
  assign _0069_ = _1241_ | _0706_;
  assign _1681_ = _1242_ | _0709_;
  assign _1683_ = _1243_ | _0712_;
  assign _1685_ = _1244_ | _0715_;
  assign _1141_[2] = _1245_ | _0718_;
  assign _0258_ = ~ { _1719_, _1719_, _1719_, _1719_ };
  assign _0259_ = ~ { _1760_, _1760_, _1760_, _1760_ };
  assign _0260_ = ~ { _1098_, _1098_, _1098_, _1098_ };
  assign _0261_ = ~ { _1762_, _1762_, _1762_, _1762_ };
  assign _0262_ = ~ { _1766_, _1766_, _1766_, _1766_ };
  assign _0263_ = ~ { _1764_, _1764_, _1764_, _1764_ };
  assign _0264_ = ~ { _1100_, _1100_, _1100_, _1100_ };
  assign _0265_ = ~ { _0426_, _0426_, _0426_, _0426_ };
  assign _0267_ = ~ _1102_;
  assign _0268_ = ~ { _1719_, _1719_, _1719_ };
  assign _0269_ = ~ { _1760_, _1760_, _1760_ };
  assign _0270_ = ~ { _1098_, _1098_, _1098_ };
  assign _0255_ = ~ _0228_;
  assign _0271_ = ~ _1104_;
  assign _0272_ = ~ _1758_;
  assign _0273_ = ~ _1106_;
  assign _0256_ = ~ _1756_;
  assign _0266_ = ~ _1759_;
  assign _0274_ = ~ { _1759_, _1759_, _1759_, _1759_, _1759_, _1759_ };
  assign _0275_ = ~ { _1719_, _1719_, _1719_, _1719_, _1719_, _1719_ };
  assign _0276_ = ~ { _0219_, _0219_ };
  assign _0277_ = ~ { _1719_, _1719_ };
  assign _0249_ = ~ _1763_;
  assign _0250_ = ~ _1762_;
  assign _0307_ = ~ ebrk_insn;
  assign _0306_ = ~ ecall_insn;
  assign _0337_ = ~ illegal_insn_q;
  assign _0311_ = ~ instr_fetch_err;
  assign _0297_ = ~ load_err_q;
  assign _0295_ = ~ store_err_q;
  assign _0338_ = ~ { _1663_, _1663_, _1663_, _1663_ };
  assign _0339_ = ~ { _1659_, _1659_, _1659_, _1659_ };
  assign _0340_ = ~ { wfi_insn, wfi_insn, wfi_insn, wfi_insn };
  assign _0316_ = ~ dret_insn;
  assign _0341_ = ~ { dret_insn, dret_insn, dret_insn };
  assign _0342_ = ~ { dret_insn, dret_insn, dret_insn, dret_insn };
  assign _0343_ = ~ { mret_insn, mret_insn, mret_insn };
  assign _0344_ = ~ { mret_insn, mret_insn, mret_insn, mret_insn };
  assign _0300_ = ~ mret_insn;
  assign _0345_ = ~ { _0416_, _0416_, _0416_, _0416_ };
  assign _0346_ = ~ _0416_;
  assign _0347_ = ~ { _0416_, _0416_, _0416_, _0416_, _0416_, _0416_ };
  assign _0348_ = ~ { load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio };
  assign _0349_ = ~ { store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio };
  assign _0350_ = ~ { ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio };
  assign _0351_ = ~ { ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio };
  assign _0352_ = ~ { illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio };
  assign _0353_ = ~ { instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio };
  assign _0354_ = ~ { load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio };
  assign _0355_ = ~ { store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio };
  assign _0356_ = ~ { ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio };
  assign _0357_ = ~ { ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio };
  assign _0358_ = ~ { illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio };
  assign _0359_ = ~ { instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio };
  assign _0360_ = ~ { ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio };
  assign _0361_ = ~ { ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio };
  assign _0362_ = ~ { illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio };
  assign _0363_ = ~ { instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio };
  assign _0364_ = ~ illegal_insn_prio;
  assign _0365_ = ~ instr_fetch_err_prio;
  assign _0366_ = ~ ebrk_insn_prio;
  assign _0367_ = ~ ecall_insn_prio;
  assign _0368_ = ~ { _1686_, _1686_, _1686_, _1686_ };
  assign _0370_ = ~ { _1686_, _1686_, _1686_, _1686_, _1686_, _1686_, _1686_, _1686_, _1686_, _1686_, _1686_, _1686_, _1686_, _1686_, _1686_, _1686_, _1686_, _1686_, _1686_, _1686_, _1686_, _1686_, _1686_, _1686_, _1686_, _1686_, _1686_, _1686_, _1686_, _1686_, _1686_, _1686_ };
  assign _0371_ = ~ { _1686_, _1686_, _1686_, _1686_, _1686_, _1686_ };
  assign _0372_ = ~ { _1686_, _1686_ };
  assign _0373_ = ~ { _1686_, _1686_, _1686_ };
  assign _0369_ = ~ _1686_;
  assign _0374_ = ~ { debug_single_step_i, debug_single_step_i, debug_single_step_i };
  assign _0375_ = ~ { trigger_match_i, trigger_match_i, trigger_match_i };
  assign _0376_ = ~ { irqs_i[17], irqs_i[17], irqs_i[17], irqs_i[17], irqs_i[17], irqs_i[17] };
  assign _0377_ = ~ { irqs_i[15], irqs_i[15], irqs_i[15], irqs_i[15], irqs_i[15], irqs_i[15] };
  assign _0378_ = ~ { _1689_, _1689_, _1689_, _1689_, _1689_, _1689_ };
  assign _0379_ = ~ { _1657_, _1657_, _1657_, _1657_, _1657_, _1657_ };
  assign _0380_ = ~ { handle_irq, handle_irq, handle_irq, handle_irq, handle_irq, handle_irq };
  assign _0291_ = ~ handle_irq;
  assign _0383_ = ~ _1655_;
  assign _0384_ = ~ { _1655_, _1655_, _1655_, _1655_ };
  assign _0385_ = ~ { _1717_, _1717_, _1717_, _1717_ };
  assign _0386_ = ~ { special_req, special_req, special_req, special_req };
  assign _0290_ = ~ enter_debug_mode;
  assign _0382_ = ~ { enter_debug_mode, enter_debug_mode, enter_debug_mode, enter_debug_mode };
  assign _0381_ = ~ { handle_irq, handle_irq, handle_irq, handle_irq };
  assign _0387_ = ~ { id_in_ready_o, id_in_ready_o, id_in_ready_o, id_in_ready_o };
  assign _0388_ = ~ { _1677_, _1677_, _1677_, _1677_ };
  assign _0254_ = ~ _1760_;
  assign _0389_ = ~ { _1758_, _1758_, _1758_ };
  assign _0390_ = ~ { _1719_, _1719_, _1719_, _1719_, _1719_, _1719_, _1719_, _1719_, _1719_, _1719_, _1719_, _1719_, _1719_, _1719_, _1719_, _1719_, _1719_, _1719_, _1719_, _1719_, _1719_, _1719_, _1719_, _1719_, _1719_, _1719_, _1719_, _1719_, _1719_, _1719_, _1719_, _1719_ };
  assign _0252_ = ~ _1719_;
  assign _0391_ = ~ { irqs_i[1], irqs_i[1], irqs_i[1], irqs_i[1] };
  assign _0392_ = ~ { irqs_i[2], irqs_i[2], irqs_i[2], irqs_i[2] };
  assign _0393_ = ~ { irqs_i[3], irqs_i[3], irqs_i[3], irqs_i[3] };
  assign _0394_ = ~ { irqs_i[4], irqs_i[4], irqs_i[4], irqs_i[4] };
  assign _0395_ = ~ { irqs_i[5], irqs_i[5], irqs_i[5], irqs_i[5] };
  assign _0396_ = ~ { irqs_i[6], irqs_i[6], irqs_i[6], irqs_i[6] };
  assign _0397_ = ~ { irqs_i[7], irqs_i[7], irqs_i[7], irqs_i[7] };
  assign _0398_ = ~ { irqs_i[8], irqs_i[8], irqs_i[8], irqs_i[8] };
  assign _0399_ = ~ { irqs_i[9], irqs_i[9], irqs_i[9], irqs_i[9] };
  assign _0400_ = ~ { irqs_i[10], irqs_i[10], irqs_i[10], irqs_i[10] };
  assign _0401_ = ~ { irqs_i[11], irqs_i[11], irqs_i[11], irqs_i[11] };
  assign _0402_ = ~ { irqs_i[12], irqs_i[12], irqs_i[12], irqs_i[12] };
  assign _0403_ = ~ { irqs_i[13], irqs_i[13], irqs_i[13], irqs_i[13] };
  assign _0404_ = ~ { irqs_i[14], irqs_i[14], irqs_i[14], irqs_i[14] };
  assign _0323_ = ~ instr_valid_i;
  assign _0405_ = ~ _1648_;
  assign _0406_ = ~ { debug_mode_o, debug_mode_o };
  assign _0407_ = ~ { instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i };
  assign _0408_ = ~ { instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i };
  assign _0409_ = ~ { _1648_, _1648_, _1648_, _1648_, _1648_, _1648_ };
  assign _1154_ = { _1141_[3], _1141_[3], _1141_[3], _1141_[3] } | _0258_;
  assign _1157_ = { controller_run_o_t0, controller_run_o_t0, controller_run_o_t0, controller_run_o_t0 } | _0259_;
  assign _1160_ = { _1099_, _1099_, _1099_, _1099_ } | _0260_;
  assign _1163_ = { _1145_[1], _1145_[1], _1145_[1], _1145_[1] } | _0261_;
  assign _1166_ = { _1767_, _1767_, _1767_, _1767_ } | _0262_;
  assign _1169_ = { _1765_, _1765_, _1765_, _1765_ } | _0263_;
  assign _1172_ = { _1101_, _1101_, _1101_, _1101_ } | _0264_;
  assign _1175_ = { _0427_, _0427_, _0427_, _0427_ } | _0265_;
  assign _1182_ = _1103_ | _0267_;
  assign _1189_ = { _1141_[3], _1141_[3], _1141_[3] } | _0268_;
  assign _1192_ = { controller_run_o_t0, controller_run_o_t0, controller_run_o_t0 } | _0269_;
  assign _1195_ = { _1099_, _1099_, _1099_ } | _0270_;
  assign _1198_ = _0229_ | _0255_;
  assign _1200_ = _1105_ | _0271_;
  assign _1204_ = _0630_ | _0272_;
  assign _1209_ = _1107_ | _0273_;
  assign _1205_ = _1757_ | _0256_;
  assign _1179_ = _1142_[1] | _0266_;
  assign _1213_ = { _1142_[1], _1142_[1], _1142_[1], _1142_[1], _1142_[1], _1142_[1] } | _0274_;
  assign _1216_ = { _1141_[3], _1141_[3], _1141_[3], _1141_[3], _1141_[3], _1141_[3] } | _0275_;
  assign _1219_ = { _0220_, _0220_ } | _0276_;
  assign _1222_ = { _1141_[3], _1141_[3] } | _0277_;
  assign _1225_ = _1145_[1] | _0250_;
  assign _1270_ = ecall_insn_t0 | _0306_;
  assign _1271_ = illegal_insn_q_t0 | _0337_;
  assign _1272_ = instr_fetch_err_t0 | _0311_;
  assign _1273_ = load_err_q_t0 | _0297_;
  assign _1274_ = store_err_prio_t0 | _0295_;
  assign _1275_ = { _1664_, _1664_, _1664_, _1664_ } | _0338_;
  assign _1278_ = { _1660_, _1660_, _1660_, _1660_ } | _0339_;
  assign _1281_ = { wfi_insn_t0, wfi_insn_t0, wfi_insn_t0, wfi_insn_t0 } | _0340_;
  assign _1284_ = { dret_insn_t0, dret_insn_t0, dret_insn_t0 } | _0341_;
  assign _1287_ = { dret_insn_t0, dret_insn_t0, dret_insn_t0, dret_insn_t0 } | _0342_;
  assign _1291_ = { mret_insn_t0, mret_insn_t0, mret_insn_t0 } | _0343_;
  assign _1294_ = { mret_insn_t0, mret_insn_t0, mret_insn_t0, mret_insn_t0 } | _0344_;
  assign _1290_ = mret_insn_t0 | _0300_;
  assign _1297_ = { _0121_, _0121_, _0121_, _0121_ } | _0345_;
  assign _1300_ = _0121_ | _0346_;
  assign _1301_ = { _0121_, _0121_, _0121_, _0121_, _0121_, _0121_ } | _0347_;
  assign _1304_ = { load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0 } | _0348_;
  assign _1307_ = { store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0 } | _0349_;
  assign _1310_ = { ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0 } | _0350_;
  assign _1313_ = { ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0 } | _0351_;
  assign _1316_ = { illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0 } | _0352_;
  assign _1319_ = { instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0 } | _0353_;
  assign _1322_ = { load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0 } | _0354_;
  assign _1325_ = { store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0 } | _0355_;
  assign _1328_ = { ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0 } | _0356_;
  assign _1331_ = { ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0 } | _0357_;
  assign _1334_ = { illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0 } | _0358_;
  assign _1337_ = { instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0 } | _0359_;
  assign _1340_ = { ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0 } | _0360_;
  assign _1343_ = { ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0 } | _0361_;
  assign _1346_ = { illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0 } | _0362_;
  assign _1349_ = { instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0 } | _0363_;
  assign _1352_ = illegal_insn_prio_t0 | _0364_;
  assign _1354_ = instr_fetch_err_prio_t0 | _0365_;
  assign _1356_ = ebrk_insn_prio_t0 | _0366_;
  assign _1359_ = ecall_insn_prio_t0 | _0367_;
  assign _1364_ = { _1141_[2], _1141_[2], _1141_[2], _1141_[2] } | _0368_;
  assign _1369_ = { _1141_[2], _1141_[2], _1141_[2], _1141_[2], _1141_[2], _1141_[2], _1141_[2], _1141_[2], _1141_[2], _1141_[2], _1141_[2], _1141_[2], _1141_[2], _1141_[2], _1141_[2], _1141_[2], _1141_[2], _1141_[2], _1141_[2], _1141_[2], _1141_[2], _1141_[2], _1141_[2], _1141_[2], _1141_[2], _1141_[2], _1141_[2], _1141_[2], _1141_[2], _1141_[2], _1141_[2], _1141_[2] } | _0370_;
  assign _1372_ = { _1141_[2], _1141_[2], _1141_[2], _1141_[2], _1141_[2], _1141_[2] } | _0371_;
  assign _1376_ = { _1141_[2], _1141_[2] } | _0372_;
  assign _1379_ = { _1141_[2], _1141_[2], _1141_[2] } | _0373_;
  assign _1367_ = _1141_[2] | _0369_;
  assign _1382_ = { debug_single_step_i_t0, debug_single_step_i_t0, debug_single_step_i_t0 } | _0374_;
  assign _1385_ = { trigger_match_i_t0, trigger_match_i_t0, trigger_match_i_t0 } | _0375_;
  assign _1388_ = { irqs_i_t0[17], irqs_i_t0[17], irqs_i_t0[17], irqs_i_t0[17], irqs_i_t0[17], irqs_i_t0[17] } | _0376_;
  assign _1391_ = { irqs_i_t0[15], irqs_i_t0[15], irqs_i_t0[15], irqs_i_t0[15], irqs_i_t0[15], irqs_i_t0[15] } | _0377_;
  assign _1394_ = { _1690_, _1690_, _1690_, _1690_, _1690_, _1690_ } | _0378_;
  assign _1397_ = { _1143_[1], _1143_[1], _1143_[1], _1143_[1], _1143_[1], _1143_[1] } | _0379_;
  assign _1401_ = { handle_irq_t0, handle_irq_t0, handle_irq_t0, handle_irq_t0, handle_irq_t0, handle_irq_t0 } | _0380_;
  assign _1400_ = handle_irq_t0 | _0291_;
  assign _1404_ = { handle_irq_t0, handle_irq_t0, handle_irq_t0, handle_irq_t0 } | _0381_;
  assign _1411_ = _1656_ | _0383_;
  assign _1414_ = { _1656_, _1656_, _1656_, _1656_ } | _0384_;
  assign _1418_ = { _1718_, _1718_, _1718_, _1718_ } | _0385_;
  assign _1421_ = { special_req_t0, special_req_t0, special_req_t0, special_req_t0 } | _0386_;
  assign _1407_ = enter_debug_mode_t0 | _0290_;
  assign _1408_ = { enter_debug_mode_t0, enter_debug_mode_t0, enter_debug_mode_t0, enter_debug_mode_t0 } | _0382_;
  assign _1426_ = { id_in_ready_o_t0, id_in_ready_o_t0, id_in_ready_o_t0, id_in_ready_o_t0 } | _0387_;
  assign _1429_ = { _0040_, _0040_, _0040_, _0040_ } | _0388_;
  assign _1432_ = { _0630_, _0630_, _0630_ } | _0389_;
  assign _1435_ = { _1141_[3], _1141_[3], _1141_[3], _1141_[3], _1141_[3], _1141_[3], _1141_[3], _1141_[3], _1141_[3], _1141_[3], _1141_[3], _1141_[3], _1141_[3], _1141_[3], _1141_[3], _1141_[3], _1141_[3], _1141_[3], _1141_[3], _1141_[3], _1141_[3], _1141_[3], _1141_[3], _1141_[3], _1141_[3], _1141_[3], _1141_[3], _1141_[3], _1141_[3], _1141_[3], _1141_[3], _1141_[3] } | _0390_;
  assign _1185_ = _1141_[3] | _0252_;
  assign _1438_ = { irqs_i_t0[1], irqs_i_t0[1], irqs_i_t0[1], irqs_i_t0[1] } | _0391_;
  assign _1441_ = { irqs_i_t0[2], irqs_i_t0[2], irqs_i_t0[2], irqs_i_t0[2] } | _0392_;
  assign _1444_ = { irqs_i_t0[3], irqs_i_t0[3], irqs_i_t0[3], irqs_i_t0[3] } | _0393_;
  assign _1447_ = { irqs_i_t0[4], irqs_i_t0[4], irqs_i_t0[4], irqs_i_t0[4] } | _0394_;
  assign _1450_ = { irqs_i_t0[5], irqs_i_t0[5], irqs_i_t0[5], irqs_i_t0[5] } | _0395_;
  assign _1453_ = { irqs_i_t0[6], irqs_i_t0[6], irqs_i_t0[6], irqs_i_t0[6] } | _0396_;
  assign _1456_ = { irqs_i_t0[7], irqs_i_t0[7], irqs_i_t0[7], irqs_i_t0[7] } | _0397_;
  assign _1459_ = { irqs_i_t0[8], irqs_i_t0[8], irqs_i_t0[8], irqs_i_t0[8] } | _0398_;
  assign _1462_ = { irqs_i_t0[9], irqs_i_t0[9], irqs_i_t0[9], irqs_i_t0[9] } | _0399_;
  assign _1465_ = { irqs_i_t0[10], irqs_i_t0[10], irqs_i_t0[10], irqs_i_t0[10] } | _0400_;
  assign _1468_ = { irqs_i_t0[11], irqs_i_t0[11], irqs_i_t0[11], irqs_i_t0[11] } | _0401_;
  assign _1471_ = { irqs_i_t0[12], irqs_i_t0[12], irqs_i_t0[12], irqs_i_t0[12] } | _0402_;
  assign _1474_ = { irqs_i_t0[13], irqs_i_t0[13], irqs_i_t0[13], irqs_i_t0[13] } | _0403_;
  assign _1477_ = { irqs_i_t0[14], irqs_i_t0[14], irqs_i_t0[14], irqs_i_t0[14] } | _0404_;
  assign _1480_ = instr_valid_i_t0 | _0323_;
  assign _1484_ = _1649_ | _0405_;
  assign _1487_ = { debug_mode_o_t0, debug_mode_o_t0 } | _0406_;
  assign _1490_ = { instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0 } | _0407_;
  assign _1493_ = { instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0 } | _0408_;
  assign _1496_ = { _1649_, _1649_, _1649_, _1649_, _1649_, _1649_ } | _0409_;
  assign _1155_ = { _1141_[3], _1141_[3], _1141_[3], _1141_[3] } | { _1719_, _1719_, _1719_, _1719_ };
  assign _1158_ = { controller_run_o_t0, controller_run_o_t0, controller_run_o_t0, controller_run_o_t0 } | { _1760_, _1760_, _1760_, _1760_ };
  assign _1161_ = { _1099_, _1099_, _1099_, _1099_ } | { _1098_, _1098_, _1098_, _1098_ };
  assign _1164_ = { _1145_[1], _1145_[1], _1145_[1], _1145_[1] } | { _1762_, _1762_, _1762_, _1762_ };
  assign _1167_ = { _1767_, _1767_, _1767_, _1767_ } | { _1766_, _1766_, _1766_, _1766_ };
  assign _1170_ = { _1765_, _1765_, _1765_, _1765_ } | { _1764_, _1764_, _1764_, _1764_ };
  assign _1173_ = { _1101_, _1101_, _1101_, _1101_ } | { _1100_, _1100_, _1100_, _1100_ };
  assign _1176_ = { _0427_, _0427_, _0427_, _0427_ } | { _0426_, _0426_, _0426_, _0426_ };
  assign _1183_ = _1103_ | _1102_;
  assign _1190_ = { _1141_[3], _1141_[3], _1141_[3] } | { _1719_, _1719_, _1719_ };
  assign _1193_ = { controller_run_o_t0, controller_run_o_t0, controller_run_o_t0 } | { _1760_, _1760_, _1760_ };
  assign _1196_ = { _1099_, _1099_, _1099_ } | { _1098_, _1098_, _1098_ };
  assign _1199_ = _1144_[3] | _1761_;
  assign _1201_ = _1105_ | _1104_;
  assign _1210_ = _1107_ | _1106_;
  assign _1206_ = _1757_ | _1756_;
  assign _1180_ = _1142_[1] | _1759_;
  assign _1214_ = { _1142_[1], _1142_[1], _1142_[1], _1142_[1], _1142_[1], _1142_[1] } | { _1759_, _1759_, _1759_, _1759_, _1759_, _1759_ };
  assign _1217_ = { _1141_[3], _1141_[3], _1141_[3], _1141_[3], _1141_[3], _1141_[3] } | { _1719_, _1719_, _1719_, _1719_, _1719_, _1719_ };
  assign _1220_ = { _0220_, _0220_ } | { _0219_, _0219_ };
  assign _1223_ = { _1141_[3], _1141_[3] } | { _1719_, _1719_ };
  assign _1226_ = _1145_[1] | _1762_;
  assign _1276_ = { _1664_, _1664_, _1664_, _1664_ } | { _1663_, _1663_, _1663_, _1663_ };
  assign _1279_ = { _1660_, _1660_, _1660_, _1660_ } | { _1659_, _1659_, _1659_, _1659_ };
  assign _1282_ = { wfi_insn_t0, wfi_insn_t0, wfi_insn_t0, wfi_insn_t0 } | { wfi_insn, wfi_insn, wfi_insn, wfi_insn };
  assign _1285_ = { dret_insn_t0, dret_insn_t0, dret_insn_t0 } | { dret_insn, dret_insn, dret_insn };
  assign _1288_ = { dret_insn_t0, dret_insn_t0, dret_insn_t0, dret_insn_t0 } | { dret_insn, dret_insn, dret_insn, dret_insn };
  assign _1292_ = { mret_insn_t0, mret_insn_t0, mret_insn_t0 } | { mret_insn, mret_insn, mret_insn };
  assign _1295_ = { mret_insn_t0, mret_insn_t0, mret_insn_t0, mret_insn_t0 } | { mret_insn, mret_insn, mret_insn, mret_insn };
  assign _1298_ = { _0121_, _0121_, _0121_, _0121_ } | { _0416_, _0416_, _0416_, _0416_ };
  assign _1302_ = { _0121_, _0121_, _0121_, _0121_, _0121_, _0121_ } | { _0416_, _0416_, _0416_, _0416_, _0416_, _0416_ };
  assign _1305_ = { load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0 } | { load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio };
  assign _1308_ = { store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0 } | { store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio };
  assign _1311_ = { ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0 } | { ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio };
  assign _1314_ = { ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0 } | { ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio };
  assign _1317_ = { illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0 } | { illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio };
  assign _1320_ = { instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0 } | { instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio };
  assign _1323_ = { load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0 } | { load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio };
  assign _1326_ = { store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0 } | { store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio };
  assign _1329_ = { ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0 } | { ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio };
  assign _1332_ = { ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0 } | { ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio };
  assign _1335_ = { illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0 } | { illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio };
  assign _1338_ = { instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0 } | { instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio };
  assign _1341_ = { ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0 } | { ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio };
  assign _1344_ = { ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0 } | { ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio };
  assign _1347_ = { illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0 } | { illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio };
  assign _1350_ = { instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0 } | { instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio };
  assign _1353_ = illegal_insn_prio_t0 | illegal_insn_prio;
  assign _1355_ = instr_fetch_err_prio_t0 | instr_fetch_err_prio;
  assign _1357_ = ebrk_insn_prio_t0 | ebrk_insn_prio;
  assign _1360_ = ecall_insn_prio_t0 | ecall_insn_prio;
  assign _1365_ = { _1141_[2], _1141_[2], _1141_[2], _1141_[2] } | { _1686_, _1686_, _1686_, _1686_ };
  assign _1370_ = { _1141_[2], _1141_[2], _1141_[2], _1141_[2], _1141_[2], _1141_[2], _1141_[2], _1141_[2], _1141_[2], _1141_[2], _1141_[2], _1141_[2], _1141_[2], _1141_[2], _1141_[2], _1141_[2], _1141_[2], _1141_[2], _1141_[2], _1141_[2], _1141_[2], _1141_[2], _1141_[2], _1141_[2], _1141_[2], _1141_[2], _1141_[2], _1141_[2], _1141_[2], _1141_[2], _1141_[2], _1141_[2] } | { _1686_, _1686_, _1686_, _1686_, _1686_, _1686_, _1686_, _1686_, _1686_, _1686_, _1686_, _1686_, _1686_, _1686_, _1686_, _1686_, _1686_, _1686_, _1686_, _1686_, _1686_, _1686_, _1686_, _1686_, _1686_, _1686_, _1686_, _1686_, _1686_, _1686_, _1686_, _1686_ };
  assign _1373_ = { _1141_[2], _1141_[2], _1141_[2], _1141_[2], _1141_[2], _1141_[2] } | { _1686_, _1686_, _1686_, _1686_, _1686_, _1686_ };
  assign _1377_ = { _1141_[2], _1141_[2] } | { _1686_, _1686_ };
  assign _1380_ = { _1141_[2], _1141_[2], _1141_[2] } | { _1686_, _1686_, _1686_ };
  assign _1368_ = _1141_[2] | _1686_;
  assign _1383_ = { debug_single_step_i_t0, debug_single_step_i_t0, debug_single_step_i_t0 } | { debug_single_step_i, debug_single_step_i, debug_single_step_i };
  assign _1386_ = { trigger_match_i_t0, trigger_match_i_t0, trigger_match_i_t0 } | { trigger_match_i, trigger_match_i, trigger_match_i };
  assign _1389_ = { irqs_i_t0[17], irqs_i_t0[17], irqs_i_t0[17], irqs_i_t0[17], irqs_i_t0[17], irqs_i_t0[17] } | { irqs_i[17], irqs_i[17], irqs_i[17], irqs_i[17], irqs_i[17], irqs_i[17] };
  assign _1392_ = { irqs_i_t0[15], irqs_i_t0[15], irqs_i_t0[15], irqs_i_t0[15], irqs_i_t0[15], irqs_i_t0[15] } | { irqs_i[15], irqs_i[15], irqs_i[15], irqs_i[15], irqs_i[15], irqs_i[15] };
  assign _1395_ = { _1690_, _1690_, _1690_, _1690_, _1690_, _1690_ } | { _1689_, _1689_, _1689_, _1689_, _1689_, _1689_ };
  assign _1398_ = { _1143_[1], _1143_[1], _1143_[1], _1143_[1], _1143_[1], _1143_[1] } | { _1657_, _1657_, _1657_, _1657_, _1657_, _1657_ };
  assign _1402_ = { handle_irq_t0, handle_irq_t0, handle_irq_t0, handle_irq_t0, handle_irq_t0, handle_irq_t0 } | { handle_irq, handle_irq, handle_irq, handle_irq, handle_irq, handle_irq };
  assign _1412_ = _1656_ | _1655_;
  assign _1415_ = { _1656_, _1656_, _1656_, _1656_ } | { _1655_, _1655_, _1655_, _1655_ };
  assign _1417_ = _0067_ | _1678_;
  assign _1419_ = { _1718_, _1718_, _1718_, _1718_ } | { _1717_, _1717_, _1717_, _1717_ };
  assign _1422_ = { special_req_t0, special_req_t0, special_req_t0, special_req_t0 } | { special_req, special_req, special_req, special_req };
  assign _1409_ = { enter_debug_mode_t0, enter_debug_mode_t0, enter_debug_mode_t0, enter_debug_mode_t0 } | { enter_debug_mode, enter_debug_mode, enter_debug_mode, enter_debug_mode };
  assign _1405_ = { handle_irq_t0, handle_irq_t0, handle_irq_t0, handle_irq_t0 } | { handle_irq, handle_irq, handle_irq, handle_irq };
  assign _1427_ = { id_in_ready_o_t0, id_in_ready_o_t0, id_in_ready_o_t0, id_in_ready_o_t0 } | { id_in_ready_o, id_in_ready_o, id_in_ready_o, id_in_ready_o };
  assign _1430_ = { _0040_, _0040_, _0040_, _0040_ } | { _1677_, _1677_, _1677_, _1677_ };
  assign _1178_ = controller_run_o_t0 | _1760_;
  assign _1433_ = { _0630_, _0630_, _0630_ } | { _1758_, _1758_, _1758_ };
  assign _1436_ = { _1141_[3], _1141_[3], _1141_[3], _1141_[3], _1141_[3], _1141_[3], _1141_[3], _1141_[3], _1141_[3], _1141_[3], _1141_[3], _1141_[3], _1141_[3], _1141_[3], _1141_[3], _1141_[3], _1141_[3], _1141_[3], _1141_[3], _1141_[3], _1141_[3], _1141_[3], _1141_[3], _1141_[3], _1141_[3], _1141_[3], _1141_[3], _1141_[3], _1141_[3], _1141_[3], _1141_[3], _1141_[3] } | { _1719_, _1719_, _1719_, _1719_, _1719_, _1719_, _1719_, _1719_, _1719_, _1719_, _1719_, _1719_, _1719_, _1719_, _1719_, _1719_, _1719_, _1719_, _1719_, _1719_, _1719_, _1719_, _1719_, _1719_, _1719_, _1719_, _1719_, _1719_, _1719_, _1719_, _1719_, _1719_ };
  assign _1186_ = _1141_[3] | _1719_;
  assign _1439_ = { irqs_i_t0[1], irqs_i_t0[1], irqs_i_t0[1], irqs_i_t0[1] } | { irqs_i[1], irqs_i[1], irqs_i[1], irqs_i[1] };
  assign _1442_ = { irqs_i_t0[2], irqs_i_t0[2], irqs_i_t0[2], irqs_i_t0[2] } | { irqs_i[2], irqs_i[2], irqs_i[2], irqs_i[2] };
  assign _1445_ = { irqs_i_t0[3], irqs_i_t0[3], irqs_i_t0[3], irqs_i_t0[3] } | { irqs_i[3], irqs_i[3], irqs_i[3], irqs_i[3] };
  assign _1448_ = { irqs_i_t0[4], irqs_i_t0[4], irqs_i_t0[4], irqs_i_t0[4] } | { irqs_i[4], irqs_i[4], irqs_i[4], irqs_i[4] };
  assign _1451_ = { irqs_i_t0[5], irqs_i_t0[5], irqs_i_t0[5], irqs_i_t0[5] } | { irqs_i[5], irqs_i[5], irqs_i[5], irqs_i[5] };
  assign _1454_ = { irqs_i_t0[6], irqs_i_t0[6], irqs_i_t0[6], irqs_i_t0[6] } | { irqs_i[6], irqs_i[6], irqs_i[6], irqs_i[6] };
  assign _1457_ = { irqs_i_t0[7], irqs_i_t0[7], irqs_i_t0[7], irqs_i_t0[7] } | { irqs_i[7], irqs_i[7], irqs_i[7], irqs_i[7] };
  assign _1460_ = { irqs_i_t0[8], irqs_i_t0[8], irqs_i_t0[8], irqs_i_t0[8] } | { irqs_i[8], irqs_i[8], irqs_i[8], irqs_i[8] };
  assign _1463_ = { irqs_i_t0[9], irqs_i_t0[9], irqs_i_t0[9], irqs_i_t0[9] } | { irqs_i[9], irqs_i[9], irqs_i[9], irqs_i[9] };
  assign _1466_ = { irqs_i_t0[10], irqs_i_t0[10], irqs_i_t0[10], irqs_i_t0[10] } | { irqs_i[10], irqs_i[10], irqs_i[10], irqs_i[10] };
  assign _1469_ = { irqs_i_t0[11], irqs_i_t0[11], irqs_i_t0[11], irqs_i_t0[11] } | { irqs_i[11], irqs_i[11], irqs_i[11], irqs_i[11] };
  assign _1472_ = { irqs_i_t0[12], irqs_i_t0[12], irqs_i_t0[12], irqs_i_t0[12] } | { irqs_i[12], irqs_i[12], irqs_i[12], irqs_i[12] };
  assign _1475_ = { irqs_i_t0[13], irqs_i_t0[13], irqs_i_t0[13], irqs_i_t0[13] } | { irqs_i[13], irqs_i[13], irqs_i[13], irqs_i[13] };
  assign _1478_ = { irqs_i_t0[14], irqs_i_t0[14], irqs_i_t0[14], irqs_i_t0[14] } | { irqs_i[14], irqs_i[14], irqs_i[14], irqs_i[14] };
  assign _1481_ = instr_valid_i_t0 | instr_valid_i;
  assign _1483_ = _1651_ | _1650_;
  assign _1485_ = _1649_ | _1648_;
  assign _1488_ = { debug_mode_o_t0, debug_mode_o_t0 } | { debug_mode_o, debug_mode_o };
  assign _1491_ = { instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0 } | { instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i };
  assign _1494_ = { instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0 } | { instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i };
  assign _1497_ = { _1649_, _1649_, _1649_, _1649_, _1649_, _1649_ } | { _1648_, _1648_, _1648_, _1648_, _1648_, _1648_ };
  assign _0571_ = 4'h0 & _1154_;
  assign _0574_ = _0135_ & _1157_;
  assign _0577_ = _1606_ & _1160_;
  assign _0580_ = 4'h0 & _1163_;
  assign _0583_ = 4'h0 & _1166_;
  assign _0586_ = _1612_ & _1169_;
  assign _0589_ = _1614_ & _1172_;
  assign _0592_ = _1616_ & _1175_;
  assign _0597_ = _1620_ & _1179_;
  assign _0600_ = _1622_ & _1182_;
  assign _0607_ = _1624_ & _1179_;
  assign _0609_ = _1626_ & _1182_;
  assign _0611_ = 3'h0 & _1189_;
  assign _0614_ = 3'h0 & _1192_;
  assign _0617_ = _1630_ & _1195_;
  assign _0620_ = _0142_ & _1198_;
  assign _0624_ = _1634_ & _1200_;
  assign _0627_ = _0224_ & _1185_;
  assign _0631_ = _0630_ & _1205_;
  assign _0634_ = _0036_ & _1185_;
  assign _0637_ = _1640_ & _1204_;
  assign _0639_ = csr_save_if_o_t0 & _1209_;
  assign _0643_ = _1642_ & _1185_;
  assign _0647_ = 6'h00 & _1213_;
  assign _0650_ = _1644_ & _1216_;
  assign _0653_ = 2'h0 & _1219_;
  assign _0656_ = _1646_ & _1222_;
  assign _0660_ = _0659_ & _1225_;
  assign _0793_ = ebrk_insn_t0 & _1270_;
  assign _0795_ = _0137_ & _1271_;
  assign _0797_ = ecall_insn_t0 & _1271_;
  assign _0799_ = _0115_ & _1272_;
  assign _0801_ = _0117_ & _1272_;
  assign _0803_ = illegal_insn_q_t0 & _1272_;
  assign _0805_ = _0090_ & _1273_;
  assign _0807_ = _0092_ & _1273_;
  assign _0809_ = _0100_ & _1273_;
  assign _0811_ = instr_fetch_err_t0 & _1273_;
  assign _0813_ = load_err_q_t0 & _1274_;
  assign _0815_ = _0047_ & _1274_;
  assign _0817_ = _0049_ & _1274_;
  assign _0819_ = _0057_ & _1274_;
  assign _0821_ = _0059_ & _1274_;
  assign _0823_ = _0005_ & _1275_;
  assign _0826_ = 4'h0 & _1278_;
  assign _0829_ = _0025_ & _1281_;
  assign _0832_ = 3'h0 & _1284_;
  assign _0835_ = _0023_ & _1287_;
  assign _0840_ = _0129_ & _1291_;
  assign _0843_ = _0021_ & _1294_;
  assign _0838_ = dret_insn_t0 & _1290_;
  assign _0847_ = 4'h0 & _1297_;
  assign _0850_ = _0083_ & _1300_;
  assign _0852_ = 6'h00 & _1301_;
  assign _0855_ = 32'd0 & _1304_;
  assign _0858_ = _1721_ & _1307_;
  assign _0861_ = _1722_ & _1310_;
  assign _0864_ = _1723_ & _1313_;
  assign _0867_ = _1725_ & _1316_;
  assign _0870_ = _1727_ & _1319_;
  assign _0873_ = 6'h00 & _1322_;
  assign _0876_ = _1729_ & _1325_;
  assign _0879_ = _1731_ & _1328_;
  assign _0882_ = _1733_ & _1331_;
  assign _0885_ = _1735_ & _1334_;
  assign _0888_ = _1737_ & _1337_;
  assign _0891_ = 4'h0 & _1340_;
  assign _0894_ = _1739_ & _1343_;
  assign _0897_ = _1741_ & _1346_;
  assign _0900_ = _1743_ & _1349_;
  assign _0903_ = _1747_ & _1352_;
  assign _0905_ = _1749_ & _1354_;
  assign _0907_ = _0083_ & _1356_;
  assign _0910_ = _1751_ & _1359_;
  assign _0913_ = _1753_ & _1352_;
  assign _0916_ = _1755_ & _1354_;
  assign _0921_ = _1745_ & _1359_;
  assign _0923_ = _0017_ & _1364_;
  assign _0928_ = 32'd0 & _1369_;
  assign _0934_ = 6'h00 & _1372_;
  assign _0937_ = _0166_ & _1367_;
  assign _0941_ = 2'h0 & _1376_;
  assign _0944_ = _0106_ & _1379_;
  assign _0947_ = _0078_ & _1367_;
  assign _0949_ = mret_insn_t0 & _1367_;
  assign _0951_ = 3'h0 & _1382_;
  assign _0954_ = _0087_ & _1385_;
  assign _0957_ = 6'h00 & _1388_;
  assign _0960_ = _0152_ & _1391_;
  assign _0963_ = _0140_ & _1394_;
  assign _0966_ = _0119_ & _1397_;
  assign _0969_ = 6'h00 & _1401_;
  assign _0972_ = _0123_ & _1400_;
  assign _0974_ = _0149_ & _1404_;
  assign _0977_ = _0162_ & _1407_;
  assign _0979_ = _0001_ & _1408_;
  assign _0982_ = _0123_ & _1411_;
  assign _0985_ = _0149_ & _1414_;
  assign _0992_ = ctrl_fsm_cs_t0 & _1418_;
  assign _0995_ = ctrl_fsm_cs_t0 & _1421_;
  assign _0998_ = handle_irq_t0 & _1407_;
  assign _1000_ = _0112_ & _1408_;
  assign _1002_ = _0085_ & _1404_;
  assign _1004_ = 4'h0 & _1426_;
  assign _1007_ = 4'h0 & _1429_;
  assign _1019_ = 3'h0 & _1432_;
  assign _1022_ = 32'd0 & _1435_;
  assign _1036_ = 4'h0 & _1438_;
  assign _1039_ = _0019_ & _1441_;
  assign _1042_ = _0015_ & _1444_;
  assign _1045_ = _0011_ & _1447_;
  assign _1048_ = _0007_ & _1450_;
  assign _1051_ = _0003_ & _1453_;
  assign _1054_ = _0178_ & _1456_;
  assign _1057_ = _0172_ & _1459_;
  assign _1060_ = _0164_ & _1462_;
  assign _1063_ = _0156_ & _1465_;
  assign _1066_ = _0144_ & _1468_;
  assign _1069_ = _0126_ & _1471_;
  assign _1072_ = _0103_ & _1474_;
  assign _1075_ = _0062_ & _1477_;
  assign _1078_ = do_single_step_q_t0 & _1480_;
  assign _1083_ = _1769_ & _1484_;
  assign _1086_ = 2'h0 & _1487_;
  assign _1089_ = pc_id_i_t0 & _1490_;
  assign _1092_ = instr_i_t0 & _1493_;
  assign _1095_ = 6'h00 & _1496_;
  assign _0572_ = _0027_ & _1155_;
  assign _0575_ = _0168_ & _1158_;
  assign _0578_ = _1604_ & _1161_;
  assign _0581_ = _0042_ & _1164_;
  assign _0584_ = 4'h0 & _1167_;
  assign _0587_ = 4'h0 & _1170_;
  assign _0590_ = _1610_ & _1173_;
  assign _0593_ = _1608_ & _1176_;
  assign _0595_ = _0069_ & _1178_;
  assign _0603_ = _0131_ & _1186_;
  assign _0605_ = _0067_ & _1178_;
  assign _0601_ = _1618_ & _1183_;
  assign _0612_ = _0065_ & _1190_;
  assign _0615_ = 3'h0 & _1193_;
  assign _0618_ = _1628_ & _1196_;
  assign _0622_ = _0098_ & _1199_;
  assign _0625_ = _1632_ & _1201_;
  assign _0628_ = _0055_ & _1186_;
  assign _0635_ = _0109_ & _1186_;
  assign _0640_ = _1638_ & _1210_;
  assign _0632_ = _0036_ & _1206_;
  assign _0644_ = _0081_ & _1186_;
  assign _0598_ = handle_irq_t0 & _1180_;
  assign _0648_ = _0051_ & _1214_;
  assign _0651_ = _0160_ & _1217_;
  assign _0654_ = 2'h0 & _1220_;
  assign _0657_ = _0053_ & _1223_;
  assign _0661_ = _0040_ & _1226_;
  assign _0824_ = 4'h0 & _1276_;
  assign _0827_ = 4'h0 & _1279_;
  assign _0830_ = 4'h0 & _1282_;
  assign _0833_ = 3'h0 & _1285_;
  assign _0836_ = 4'h0 & _1288_;
  assign _0841_ = 3'h0 & _1292_;
  assign _0844_ = 4'h0 & _1295_;
  assign _0848_ = 4'h0 & _1298_;
  assign _0853_ = 6'h00 & _1302_;
  assign _0856_ = lsu_addr_last_i_t0 & _1305_;
  assign _0859_ = lsu_addr_last_i_t0 & _1308_;
  assign _0862_ = 32'd0 & _1311_;
  assign _0865_ = 32'd0 & _1314_;
  assign _0868_ = _1775_ & _1317_;
  assign _0871_ = _1773_ & _1320_;
  assign _0874_ = 6'h00 & _1323_;
  assign _0877_ = 6'h00 & _1326_;
  assign _0880_ = _0176_ & _1329_;
  assign _0883_ = _1777_ & _1332_;
  assign _0886_ = 6'h00 & _1335_;
  assign _0889_ = 6'h00 & _1338_;
  assign _0892_ = _0013_ & _1341_;
  assign _0895_ = 4'h0 & _1344_;
  assign _0898_ = 4'h0 & _1347_;
  assign _0901_ = 4'h0 & _1350_;
  assign _0908_ = _0147_ & _1357_;
  assign _0911_ = _0083_ & _1360_;
  assign _0914_ = _0083_ & _1353_;
  assign _0917_ = _0083_ & _1355_;
  assign _0919_ = _0121_ & _1357_;
  assign _0924_ = _0009_ & _1365_;
  assign _0929_ = _0076_ & _1370_;
  assign _0932_ = _0133_ & _1368_;
  assign _0935_ = _0170_ & _1373_;
  assign _0926_ = _0096_ & _1368_;
  assign _0939_ = _0083_ & _1368_;
  assign _0942_ = _1771_ & _1377_;
  assign _0945_ = 3'h0 & _1380_;
  assign _0952_ = 3'h0 & _1383_;
  assign _0955_ = 3'h0 & _1386_;
  assign _0958_ = 6'h00 & _1389_;
  assign _0961_ = 6'h00 & _1392_;
  assign _0964_ = { 2'h0, mfip_id_t0 } & _1395_;
  assign _0967_ = 6'h00 & _1398_;
  assign _0970_ = _0094_ & _1402_;
  assign _0983_ = _0154_ & _1412_;
  assign _0986_ = _0174_ & _1415_;
  assign _0988_ = jump_set_i_t0 & _1417_;
  assign _0990_ = branch_set_i_t0 & _1417_;
  assign _0993_ = 4'h0 & _1419_;
  assign _0996_ = _0158_ & _1422_;
  assign _0980_ = 4'h0 & _1409_;
  assign _0975_ = 4'h0 & _1405_;
  assign _1005_ = 4'h0 & _1427_;
  assign _1008_ = 4'h0 & _1430_;
  assign _1011_ = special_req_t0 & _1178_;
  assign _1014_ = _0073_ & _1178_;
  assign _1016_ = _0071_ & _1178_;
  assign _1020_ = _0044_ & _1433_;
  assign _1023_ = _0029_ & _1436_;
  assign _1025_ = _0031_ & _1186_;
  assign _1027_ = _0033_ & _1186_;
  assign _1029_ = _0038_ & _1186_;
  assign _1037_ = 4'h0 & _1439_;
  assign _1040_ = 4'h0 & _1442_;
  assign _1043_ = 4'h0 & _1445_;
  assign _1046_ = 4'h0 & _1448_;
  assign _1049_ = 4'h0 & _1451_;
  assign _1052_ = 4'h0 & _1454_;
  assign _1055_ = 4'h0 & _1457_;
  assign _1058_ = 4'h0 & _1460_;
  assign _1061_ = 4'h0 & _1463_;
  assign _1064_ = 4'h0 & _1466_;
  assign _1067_ = 4'h0 & _1469_;
  assign _1070_ = 4'h0 & _1472_;
  assign _1073_ = 4'h0 & _1475_;
  assign _1076_ = 4'h0 & _1478_;
  assign _1079_ = _0184_ & _1481_;
  assign _1081_ = debug_ebreaku_i_t0 & _1483_;
  assign _1084_ = debug_ebreakm_i_t0 & _1485_;
  assign _1087_ = 2'h0 & _1488_;
  assign _1090_ = _0180_ & _1491_;
  assign _1093_ = { 16'h0000, instr_compressed_i_t0 } & _1494_;
  assign _1096_ = 6'h00 & _1497_;
  assign _1156_ = _0571_ | _0572_;
  assign _1159_ = _0574_ | _0575_;
  assign _1162_ = _0577_ | _0578_;
  assign _1165_ = _0580_ | _0581_;
  assign _1168_ = _0583_ | _0584_;
  assign _1171_ = _0586_ | _0587_;
  assign _1174_ = _0589_ | _0590_;
  assign _1177_ = _0592_ | _0593_;
  assign _1181_ = _0597_ | _0598_;
  assign _1184_ = _0600_ | _0601_;
  assign _1187_ = _0607_ | _0598_;
  assign _1188_ = _0609_ | _0601_;
  assign _1191_ = _0611_ | _0612_;
  assign _1194_ = _0614_ | _0615_;
  assign _1197_ = _0617_ | _0618_;
  assign _1202_ = _0624_ | _0625_;
  assign _1203_ = _0627_ | _0628_;
  assign _1207_ = _0631_ | _0632_;
  assign _1208_ = _0634_ | _0635_;
  assign _1211_ = _0639_ | _0640_;
  assign _1212_ = _0643_ | _0644_;
  assign _1215_ = _0647_ | _0648_;
  assign _1218_ = _0650_ | _0651_;
  assign _1221_ = _0653_ | _0654_;
  assign _1224_ = _0656_ | _0657_;
  assign _1227_ = _0660_ | _0661_;
  assign _1277_ = _0823_ | _0824_;
  assign _1280_ = _0826_ | _0827_;
  assign _1283_ = _0829_ | _0830_;
  assign _1286_ = _0832_ | _0833_;
  assign _1289_ = _0835_ | _0836_;
  assign _1293_ = _0840_ | _0841_;
  assign _1296_ = _0843_ | _0844_;
  assign _1299_ = _0847_ | _0848_;
  assign _1303_ = _0852_ | _0853_;
  assign _1306_ = _0855_ | _0856_;
  assign _1309_ = _0858_ | _0859_;
  assign _1312_ = _0861_ | _0862_;
  assign _1315_ = _0864_ | _0865_;
  assign _1318_ = _0867_ | _0868_;
  assign _1321_ = _0870_ | _0871_;
  assign _1324_ = _0873_ | _0874_;
  assign _1327_ = _0876_ | _0877_;
  assign _1330_ = _0879_ | _0880_;
  assign _1333_ = _0882_ | _0883_;
  assign _1336_ = _0885_ | _0886_;
  assign _1339_ = _0888_ | _0889_;
  assign _1342_ = _0891_ | _0892_;
  assign _1345_ = _0894_ | _0895_;
  assign _1348_ = _0897_ | _0898_;
  assign _1351_ = _0900_ | _0901_;
  assign _1358_ = _0907_ | _0908_;
  assign _1361_ = _0910_ | _0911_;
  assign _1362_ = _0913_ | _0914_;
  assign _1363_ = _0916_ | _0917_;
  assign _1366_ = _0923_ | _0924_;
  assign _1371_ = _0928_ | _0929_;
  assign _1374_ = _0934_ | _0935_;
  assign _1375_ = _0937_ | _0926_;
  assign _1378_ = _0941_ | _0942_;
  assign _1381_ = _0944_ | _0945_;
  assign _1384_ = _0951_ | _0952_;
  assign _1387_ = _0954_ | _0955_;
  assign _1390_ = _0957_ | _0958_;
  assign _1393_ = _0960_ | _0961_;
  assign _1396_ = _0963_ | _0964_;
  assign _1399_ = _0966_ | _0967_;
  assign _1403_ = _0969_ | _0970_;
  assign _1406_ = _0974_ | _0975_;
  assign _1410_ = _0979_ | _0980_;
  assign _1413_ = _0982_ | _0983_;
  assign _1416_ = _0985_ | _0986_;
  assign _1420_ = _0992_ | _0993_;
  assign _1423_ = _0995_ | _0996_;
  assign _1424_ = _1000_ | _0980_;
  assign _1425_ = _1002_ | _0975_;
  assign _1428_ = _1004_ | _1005_;
  assign _1431_ = _1007_ | _1008_;
  assign _1434_ = _1019_ | _1020_;
  assign _1437_ = _1022_ | _1023_;
  assign _1440_ = _1036_ | _1037_;
  assign _1443_ = _1039_ | _1040_;
  assign _1446_ = _1042_ | _1043_;
  assign _1449_ = _1045_ | _1046_;
  assign _1452_ = _1048_ | _1049_;
  assign _1455_ = _1051_ | _1052_;
  assign _1458_ = _1054_ | _1055_;
  assign _1461_ = _1057_ | _1058_;
  assign _1464_ = _1060_ | _1061_;
  assign _1467_ = _1063_ | _1064_;
  assign _1470_ = _1066_ | _1067_;
  assign _1473_ = _1069_ | _1070_;
  assign _1476_ = _1072_ | _1073_;
  assign _1479_ = _1075_ | _1076_;
  assign _1482_ = _1078_ | _1079_;
  assign _1486_ = _1083_ | _1084_;
  assign _1489_ = _1086_ | _1087_;
  assign _1492_ = _1089_ | _1090_;
  assign _1495_ = _1092_ | _1093_;
  assign _1498_ = _1095_ | _1096_;
  assign _1503_ = 4'h5 ^ _0026_;
  assign _1504_ = _0134_ ^ _0167_;
  assign _1505_ = _1605_ ^ _1603_;
  assign _1506_ = 4'h3 ^ _0041_;
  assign _1507_ = _1611_ ^ 4'h4;
  assign _1508_ = _1613_ ^ _1609_;
  assign _1509_ = _1615_ ^ _1607_;
  assign _1510_ = _1619_ ^ _0034_;
  assign _1511_ = _1621_ ^ _1617_;
  assign _1512_ = _1623_ ^ _0034_;
  assign _1513_ = _1625_ ^ _1617_;
  assign _1514_ = 3'h2 ^ _0064_;
  assign _1515_ = _1629_ ^ _1627_;
  assign _1516_ = _1633_ ^ _1631_;
  assign _1517_ = _0063_ ^ _0127_;
  assign _1518_ = _1635_ ^ _0054_;
  assign _1519_ = _1636_ ^ _0035_;
  assign _1520_ = _0035_ ^ _0108_;
  assign _1521_ = csr_save_if_o ^ _1637_;
  assign _1522_ = _1641_ ^ _0080_;
  assign _1523_ = _1643_ ^ _0159_;
  assign _1524_ = _1645_ ^ _0052_;
  assign _1525_ = _1647_ ^ _0039_;
  assign _1526_ = _0004_ ^ 4'h8;
  assign _1527_ = _0024_ ^ 4'h2;
  assign _1528_ = _0022_ ^ 4'h5;
  assign _1529_ = _0128_ ^ 3'h3;
  assign _1530_ = _0020_ ^ 4'h5;
  assign _1531_ = _1720_ ^ lsu_addr_last_i;
  assign _1534_ = _1724_ ^ _1774_;
  assign _1535_ = _1726_ ^ _1772_;
  assign _1536_ = _1728_ ^ 6'h07;
  assign _1537_ = _1730_ ^ _0175_;
  assign _1538_ = _1732_ ^ _1776_;
  assign _1539_ = _1734_ ^ 6'h02;
  assign _1540_ = _1736_ ^ 6'h01;
  assign _1541_ = 4'h5 ^ _0012_;
  assign _1542_ = _1738_ ^ 4'h5;
  assign _1543_ = _1740_ ^ 4'h5;
  assign _1544_ = _1742_ ^ 4'h5;
  assign _1545_ = _0110_ ^ _0146_;
  assign _1546_ = _1750_ ^ _0110_;
  assign _1547_ = _1752_ ^ _0110_;
  assign _1548_ = _1754_ ^ _0110_;
  assign _1549_ = _0016_ ^ _0008_;
  assign _1550_ = _0165_ ^ _0095_;
  assign _1551_ = 2'h1 ^ _1770_;
  assign _1552_ = _0105_ ^ 3'h2;
  assign _1553_ = _0086_ ^ 3'h2;
  assign _1554_ = _0151_ ^ 6'h2b;
  assign _1555_ = _0139_ ^ { 2'h3, mfip_id };
  assign _1556_ = _0118_ ^ 6'h3f;
  assign _1557_ = _0148_ ^ 4'h7;
  assign _1558_ = _0000_ ^ 4'h8;
  assign _1559_ = _0122_ ^ _0153_;
  assign _1560_ = _0148_ ^ _0173_;
  assign _1561_ = ctrl_fsm_cs ^ 4'h6;
  assign _1562_ = ctrl_fsm_cs ^ _0157_;
  assign _1563_ = _0111_ ^ 4'h8;
  assign _1564_ = _0084_ ^ 4'h7;
  assign _1565_ = 3'h1 ^ _0043_;
  assign _1566_ = _0018_ ^ 4'h2;
  assign _1567_ = _0014_ ^ 4'h3;
  assign _1568_ = _0010_ ^ 4'h4;
  assign _1569_ = _0006_ ^ 4'h5;
  assign _1570_ = _0002_ ^ 4'h6;
  assign _1571_ = _0177_ ^ 4'h7;
  assign _1572_ = _0171_ ^ 4'h8;
  assign _1573_ = _0163_ ^ 4'h9;
  assign _1574_ = _0155_ ^ 4'ha;
  assign _1575_ = _0143_ ^ 4'hb;
  assign _1576_ = _0125_ ^ 4'hc;
  assign _1577_ = _0102_ ^ 4'hd;
  assign _1578_ = _0061_ ^ 4'he;
  assign _1579_ = do_single_step_q ^ _0183_;
  assign _1580_ = _1768_ ^ debug_ebreakm_i;
  assign _1581_ = pc_id_i ^ _0179_;
  assign _1582_ = instr_i ^ { 16'h0000, instr_compressed_i };
  assign _0573_ = { _1141_[3], _1141_[3], _1141_[3], _1141_[3] } & _1503_;
  assign _0576_ = { controller_run_o_t0, controller_run_o_t0, controller_run_o_t0, controller_run_o_t0 } & _1504_;
  assign _0579_ = { _1099_, _1099_, _1099_, _1099_ } & _1505_;
  assign _0582_ = { _1145_[1], _1145_[1], _1145_[1], _1145_[1] } & _1506_;
  assign _0585_ = { _1767_, _1767_, _1767_, _1767_ } & 4'h1;
  assign _0588_ = { _1765_, _1765_, _1765_, _1765_ } & _1507_;
  assign _0591_ = { _1101_, _1101_, _1101_, _1101_ } & _1508_;
  assign _0594_ = { _0427_, _0427_, _0427_, _0427_ } & _1509_;
  assign _0596_ = controller_run_o_t0 & _0068_;
  assign _0599_ = _1142_[1] & _1510_;
  assign _0602_ = _1103_ & _1511_;
  assign _0604_ = _1141_[3] & _0420_;
  assign _0606_ = controller_run_o_t0 & _0066_;
  assign _0608_ = _1142_[1] & _1512_;
  assign _0610_ = _1103_ & _1513_;
  assign _0613_ = { _1141_[3], _1141_[3], _1141_[3] } & _1514_;
  assign _0616_ = { controller_run_o_t0, controller_run_o_t0, controller_run_o_t0 } & 3'h1;
  assign _0619_ = { _1099_, _1099_, _1099_ } & _1515_;
  assign _0621_ = _0229_ & _0413_;
  assign _0623_ = _1144_[3] & _0097_;
  assign _0626_ = _1105_ & _1516_;
  assign debug_mode_d_t0 = _1141_[3] & _0414_;
  assign nmi_mode_d_t0 = _1141_[3] & _1517_;
  assign _0629_ = _1141_[3] & _1518_;
  assign _0633_ = _1757_ & _1519_;
  assign _0636_ = _1141_[3] & _1520_;
  assign _0638_ = _0630_ & _0422_;
  assign _0641_ = _1107_ & _1521_;
  assign _0642_ = _1757_ & _0035_;
  assign _0645_ = _1141_[3] & _1522_;
  assign _0646_ = _1142_[1] & _0034_;
  assign _0649_ = { _1142_[1], _1142_[1], _1142_[1], _1142_[1], _1142_[1], _1142_[1] } & _0050_;
  assign _0652_ = { _1141_[3], _1141_[3], _1141_[3], _1141_[3], _1141_[3], _1141_[3] } & _1523_;
  assign _0655_ = { _0220_, _0220_ } & 2'h3;
  assign _0658_ = { _1141_[3], _1141_[3] } & _1524_;
  assign _0662_ = _1145_[1] & _1525_;
  assign _0794_ = ecall_insn_t0 & _0150_;
  assign _0796_ = illegal_insn_q_t0 & _0136_;
  assign _0798_ = illegal_insn_q_t0 & _0138_;
  assign _0800_ = instr_fetch_err_t0 & _0114_;
  assign _0802_ = instr_fetch_err_t0 & _0116_;
  assign _0804_ = instr_fetch_err_t0 & _0124_;
  assign _0806_ = load_err_q_t0 & _0089_;
  assign _0808_ = load_err_q_t0 & _0091_;
  assign _0810_ = load_err_q_t0 & _0099_;
  assign _0812_ = load_err_q_t0 & _0101_;
  assign _0814_ = store_err_prio_t0 & _0060_;
  assign _0816_ = store_err_prio_t0 & _0046_;
  assign _0818_ = store_err_prio_t0 & _0048_;
  assign _0820_ = store_err_prio_t0 & _0056_;
  assign _0822_ = store_err_prio_t0 & _0058_;
  assign _0825_ = { _1664_, _1664_, _1664_, _1664_ } & _1526_;
  assign _0828_ = { _1660_, _1660_, _1660_, _1660_ } & 4'h2;
  assign _0831_ = { wfi_insn_t0, wfi_insn_t0, wfi_insn_t0, wfi_insn_t0 } & _1527_;
  assign _0834_ = { dret_insn_t0, dret_insn_t0, dret_insn_t0 } & 3'h4;
  assign _0837_ = { dret_insn_t0, dret_insn_t0, dret_insn_t0, dret_insn_t0 } & _1528_;
  assign _0839_ = mret_insn_t0 & _0415_;
  assign _0842_ = { mret_insn_t0, mret_insn_t0, mret_insn_t0 } & _1529_;
  assign _0845_ = { mret_insn_t0, mret_insn_t0, mret_insn_t0, mret_insn_t0 } & _1530_;
  assign _0846_ = mret_insn_t0 & _0107_;
  assign _0849_ = { _0121_, _0121_, _0121_, _0121_ } & 4'hc;
  assign _0851_ = _0121_ & _0110_;
  assign _0854_ = { _0121_, _0121_, _0121_, _0121_, _0121_, _0121_ } & 6'h03;
  assign _0857_ = { load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0 } & lsu_addr_last_i;
  assign _0860_ = { store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0 } & _1531_;
  assign _0863_ = { ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0 } & _1532_;
  assign _0866_ = { ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0 } & _1533_;
  assign _0869_ = { illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0 } & _1534_;
  assign _0872_ = { instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0 } & _1535_;
  assign _0875_ = { load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0 } & 6'h05;
  assign _0878_ = { store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0 } & _1536_;
  assign _0881_ = { ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0 } & _1537_;
  assign _0884_ = { ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0 } & _1538_;
  assign _0887_ = { illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0 } & _1539_;
  assign _0890_ = { instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0 } & _1540_;
  assign _0893_ = { ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0 } & _1541_;
  assign _0896_ = { ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0 } & _1542_;
  assign _0899_ = { illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0 } & _1543_;
  assign _0902_ = { instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0 } & _1544_;
  assign _0904_ = illegal_insn_prio_t0 & _0418_;
  assign _0906_ = instr_fetch_err_prio_t0 & _0419_;
  assign _0909_ = ebrk_insn_prio_t0 & _1545_;
  assign _0912_ = ecall_insn_prio_t0 & _1546_;
  assign _0915_ = illegal_insn_prio_t0 & _1547_;
  assign _0918_ = instr_fetch_err_prio_t0 & _1548_;
  assign _0920_ = ebrk_insn_prio_t0 & _0416_;
  assign _0922_ = ecall_insn_prio_t0 & _0417_;
  assign _0925_ = { _1141_[2], _1141_[2], _1141_[2], _1141_[2] } & _1549_;
  assign _0927_ = _1141_[2] & _0421_;
  assign _0930_ = { _1141_[2], _1141_[2], _1141_[2], _1141_[2], _1141_[2], _1141_[2], _1141_[2], _1141_[2], _1141_[2], _1141_[2], _1141_[2], _1141_[2], _1141_[2], _1141_[2], _1141_[2], _1141_[2], _1141_[2], _1141_[2], _1141_[2], _1141_[2], _1141_[2], _1141_[2], _1141_[2], _1141_[2], _1141_[2], _1141_[2], _1141_[2], _1141_[2], _1141_[2], _1141_[2], _1141_[2], _1141_[2] } & _0075_;
  assign _0931_ = _1141_[2] & _0095_;
  assign _0933_ = _1141_[2] & _0132_;
  assign _0936_ = { _1141_[2], _1141_[2], _1141_[2], _1141_[2], _1141_[2], _1141_[2] } & _0169_;
  assign _0938_ = _1141_[2] & _1550_;
  assign _0940_ = _1141_[2] & _0082_;
  assign _0943_ = { _1141_[2], _1141_[2] } & _1551_;
  assign _0946_ = { _1141_[2], _1141_[2], _1141_[2] } & _1552_;
  assign _0948_ = _1141_[2] & _0077_;
  assign _0950_ = _1141_[2] & _0079_;
  assign _0953_ = { debug_single_step_i_t0, debug_single_step_i_t0, debug_single_step_i_t0 } & 3'h7;
  assign _0956_ = { trigger_match_i_t0, trigger_match_i_t0, trigger_match_i_t0 } & _1553_;
  assign _0959_ = { irqs_i_t0[17], irqs_i_t0[17], irqs_i_t0[17], irqs_i_t0[17], irqs_i_t0[17], irqs_i_t0[17] } & 6'h04;
  assign _0962_ = { irqs_i_t0[15], irqs_i_t0[15], irqs_i_t0[15], irqs_i_t0[15], irqs_i_t0[15], irqs_i_t0[15] } & _1554_;
  assign _0965_ = { _1690_, _1690_, _1690_, _1690_, _1690_, _1690_ } & _1555_;
  assign _0968_ = { _1143_[1], _1143_[1], _1143_[1], _1143_[1], _1143_[1], _1143_[1] } & _1556_;
  assign _0971_ = { handle_irq_t0, handle_irq_t0, handle_irq_t0, handle_irq_t0, handle_irq_t0, handle_irq_t0 } & _0093_;
  assign _0973_ = handle_irq_t0 & _0411_;
  assign _0976_ = { handle_irq_t0, handle_irq_t0, handle_irq_t0, handle_irq_t0 } & _1557_;
  assign _0978_ = enter_debug_mode_t0 & _0412_;
  assign _0981_ = { enter_debug_mode_t0, enter_debug_mode_t0, enter_debug_mode_t0, enter_debug_mode_t0 } & _1558_;
  assign _0984_ = _1656_ & _1559_;
  assign _0987_ = { _1656_, _1656_, _1656_, _1656_ } & _1560_;
  assign _0989_ = _0067_ & jump_set_i;
  assign _0991_ = _0067_ & branch_set_i;
  assign _0994_ = { _1718_, _1718_, _1718_, _1718_ } & _1561_;
  assign _0997_ = { special_req_t0, special_req_t0, special_req_t0, special_req_t0 } & _1562_;
  assign _0999_ = enter_debug_mode_t0 & _0410_;
  assign _1001_ = { enter_debug_mode_t0, enter_debug_mode_t0, enter_debug_mode_t0, enter_debug_mode_t0 } & _1563_;
  assign _1003_ = { handle_irq_t0, handle_irq_t0, handle_irq_t0, handle_irq_t0 } & _1564_;
  assign _1006_ = { id_in_ready_o_t0, id_in_ready_o_t0, id_in_ready_o_t0, id_in_ready_o_t0 } & 4'hx;
  assign _1009_ = { _0040_, _0040_, _0040_, _0040_ } & 4'hx;
  assign _1012_ = controller_run_o_t0 & _0074_;
  assign _1015_ = controller_run_o_t0 & _0072_;
  assign _1017_ = controller_run_o_t0 & _0070_;
  assign _1021_ = { _0630_, _0630_, _0630_ } & _1565_;
  assign _1024_ = { _1141_[3], _1141_[3], _1141_[3], _1141_[3], _1141_[3], _1141_[3], _1141_[3], _1141_[3], _1141_[3], _1141_[3], _1141_[3], _1141_[3], _1141_[3], _1141_[3], _1141_[3], _1141_[3], _1141_[3], _1141_[3], _1141_[3], _1141_[3], _1141_[3], _1141_[3], _1141_[3], _1141_[3], _1141_[3], _1141_[3], _1141_[3], _1141_[3], _1141_[3], _1141_[3], _1141_[3], _1141_[3] } & _0028_;
  assign _1026_ = _1141_[3] & _0030_;
  assign _1028_ = _1141_[3] & _0032_;
  assign _1030_ = _1141_[3] & _0037_;
  assign _1038_ = { irqs_i_t0[1], irqs_i_t0[1], irqs_i_t0[1], irqs_i_t0[1] } & 4'h1;
  assign _1041_ = { irqs_i_t0[2], irqs_i_t0[2], irqs_i_t0[2], irqs_i_t0[2] } & _1566_;
  assign _1044_ = { irqs_i_t0[3], irqs_i_t0[3], irqs_i_t0[3], irqs_i_t0[3] } & _1567_;
  assign _1047_ = { irqs_i_t0[4], irqs_i_t0[4], irqs_i_t0[4], irqs_i_t0[4] } & _1568_;
  assign _1050_ = { irqs_i_t0[5], irqs_i_t0[5], irqs_i_t0[5], irqs_i_t0[5] } & _1569_;
  assign _1053_ = { irqs_i_t0[6], irqs_i_t0[6], irqs_i_t0[6], irqs_i_t0[6] } & _1570_;
  assign _1056_ = { irqs_i_t0[7], irqs_i_t0[7], irqs_i_t0[7], irqs_i_t0[7] } & _1571_;
  assign _1059_ = { irqs_i_t0[8], irqs_i_t0[8], irqs_i_t0[8], irqs_i_t0[8] } & _1572_;
  assign _1062_ = { irqs_i_t0[9], irqs_i_t0[9], irqs_i_t0[9], irqs_i_t0[9] } & _1573_;
  assign _1065_ = { irqs_i_t0[10], irqs_i_t0[10], irqs_i_t0[10], irqs_i_t0[10] } & _1574_;
  assign _1068_ = { irqs_i_t0[11], irqs_i_t0[11], irqs_i_t0[11], irqs_i_t0[11] } & _1575_;
  assign _1071_ = { irqs_i_t0[12], irqs_i_t0[12], irqs_i_t0[12], irqs_i_t0[12] } & _1576_;
  assign _1074_ = { irqs_i_t0[13], irqs_i_t0[13], irqs_i_t0[13], irqs_i_t0[13] } & _1577_;
  assign _1077_ = { irqs_i_t0[14], irqs_i_t0[14], irqs_i_t0[14], irqs_i_t0[14] } & _1578_;
  assign _1080_ = instr_valid_i_t0 & _1579_;
  assign _1082_ = _1651_ & debug_ebreaku_i;
  assign _1085_ = _1649_ & _1580_;
  assign _1088_ = { debug_mode_o_t0, debug_mode_o_t0 } & 2'h3;
  assign _1091_ = { instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0 } & _1581_;
  assign _1094_ = { instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0 } & _1582_;
  assign _1097_ = { _1649_, _1649_, _1649_, _1649_, _1649_, _1649_ } & 6'h03;
  assign _1604_ = _0573_ | _1156_;
  assign _1606_ = _0576_ | _1159_;
  assign _1608_ = _0579_ | _1162_;
  assign _1610_ = _0582_ | _1165_;
  assign _1612_ = _0585_ | _1168_;
  assign _1614_ = _0588_ | _1171_;
  assign _1616_ = _0591_ | _1174_;
  assign ctrl_fsm_ns_t0 = _0594_ | _1177_;
  assign _1620_ = _0596_ | _0595_;
  assign _1622_ = _0599_ | _1181_;
  assign pc_set_spec_o_t0 = _0602_ | _1184_;
  assign _1618_ = _0604_ | _0603_;
  assign _1624_ = _0606_ | _0605_;
  assign _1626_ = _0608_ | _1187_;
  assign pc_set_o_t0 = _0610_ | _1188_;
  assign _1628_ = _0613_ | _1191_;
  assign _1630_ = _0616_ | _1194_;
  assign pc_mux_o_t0 = _0619_ | _1197_;
  assign _1632_ = _0621_ | _0620_;
  assign _1634_ = _0623_ | _0622_;
  assign halt_if_t0 = _0626_ | _1202_;
  assign flush_id_o_t0 = _0629_ | _1203_;
  assign debug_csr_save_o_t0 = _0633_ | _1207_;
  assign _1638_ = _0636_ | _1208_;
  assign csr_save_if_o_t0 = _0638_ | _0637_;
  assign csr_save_cause_o_t0 = _0641_ | _1211_;
  assign _1642_ = _0642_ | _0632_;
  assign csr_save_id_o_t0 = _0645_ | _1212_;
  assign _1640_ = _0646_ | _0598_;
  assign _1644_ = _0649_ | _1215_;
  assign exc_cause_o_t0 = _0652_ | _1218_;
  assign _1646_ = _0655_ | _1221_;
  assign exc_pc_mux_o_t0 = _0658_ | _1224_;
  assign ctrl_busy_o_t0 = _0662_ | _1227_;
  assign _0137_ = _0794_ | _0793_;
  assign _0115_ = _0796_ | _0795_;
  assign _0117_ = _0798_ | _0797_;
  assign _0090_ = _0800_ | _0799_;
  assign _0092_ = _0802_ | _0801_;
  assign _0100_ = _0804_ | _0803_;
  assign _0047_ = _0806_ | _0805_;
  assign _0049_ = _0808_ | _0807_;
  assign _0057_ = _0810_ | _0809_;
  assign _0059_ = _0812_ | _0811_;
  assign load_err_prio_t0 = _0814_ | _0813_;
  assign ebrk_insn_prio_t0 = _0816_ | _0815_;
  assign ecall_insn_prio_t0 = _0818_ | _0817_;
  assign illegal_insn_prio_t0 = _0820_ | _0819_;
  assign instr_fetch_err_prio_t0 = _0822_ | _0821_;
  assign _0027_ = _0825_ | _1277_;
  assign _0025_ = _0828_ | _1280_;
  assign _0023_ = _0831_ | _1283_;
  assign _0129_ = _0834_ | _1286_;
  assign _0021_ = _0837_ | _1289_;
  assign _0166_ = _0839_ | _0838_;
  assign _0106_ = _0842_ | _1293_;
  assign _0017_ = _0845_ | _1296_;
  assign _0078_ = _0846_ | _0838_;
  assign _0013_ = _0849_ | _1299_;
  assign _0147_ = _0851_ | _0850_;
  assign _0176_ = _0854_ | _1303_;
  assign _1721_ = _0857_ | _1306_;
  assign _1722_ = _0860_ | _1309_;
  assign _1723_ = _0863_ | _1312_;
  assign _1725_ = _0866_ | _1315_;
  assign _1727_ = _0869_ | _1318_;
  assign _0076_ = _0872_ | _1321_;
  assign _1729_ = _0875_ | _1324_;
  assign _1731_ = _0878_ | _1327_;
  assign _1733_ = _0881_ | _1330_;
  assign _1735_ = _0884_ | _1333_;
  assign _1737_ = _0887_ | _1336_;
  assign _0170_ = _0890_ | _1339_;
  assign _1739_ = _0893_ | _1342_;
  assign _1741_ = _0896_ | _1345_;
  assign _1743_ = _0899_ | _1348_;
  assign _0009_ = _0902_ | _1351_;
  assign _1749_ = _0904_ | _0903_;
  assign _0096_ = _0906_ | _0905_;
  assign _1751_ = _0909_ | _1358_;
  assign _1753_ = _0912_ | _1361_;
  assign _1755_ = _0915_ | _1362_;
  assign _0133_ = _0918_ | _1363_;
  assign _1745_ = _0920_ | _0919_;
  assign _1747_ = _0922_ | _0921_;
  assign _0005_ = _0925_ | _1366_;
  assign _0055_ = _0927_ | _0926_;
  assign _0029_ = _0930_ | _1371_;
  assign _0109_ = _0931_ | _0926_;
  assign _0081_ = _0933_ | _0932_;
  assign _0160_ = _0936_ | _1374_;
  assign _0131_ = _0938_ | _1375_;
  assign _0038_ = _0940_ | _0939_;
  assign _0053_ = _0943_ | _1378_;
  assign _0065_ = _0946_ | _1381_;
  assign _0031_ = _0948_ | _0947_;
  assign _0033_ = _0950_ | _0949_;
  assign _0087_ = _0953_ | _1384_;
  assign _0044_ = _0956_ | _1387_;
  assign _0152_ = _0959_ | _1390_;
  assign _0140_ = _0962_ | _1393_;
  assign _0119_ = _0965_ | _1396_;
  assign _0094_ = _0968_ | _1399_;
  assign _0051_ = _0971_ | _1403_;
  assign _0162_ = _0973_ | _0972_;
  assign _0001_ = _0976_ | _1406_;
  assign _0154_ = _0978_ | _0977_;
  assign _0174_ = _0981_ | _1410_;
  assign _0142_ = _0984_ | _1413_;
  assign _0168_ = _0987_ | _1416_;
  assign _0071_ = _0989_ | _0988_;
  assign _0073_ = _0991_ | _0990_;
  assign _0158_ = _0994_ | _1420_;
  assign _0149_ = _0997_ | _1423_;
  assign _0098_ = _0999_ | _0998_;
  assign _0135_ = _1001_ | _1424_;
  assign _0112_ = _1003_ | _1425_;
  assign _0085_ = _1006_ | _1428_;
  assign _0042_ = _1009_ | _1431_;
  assign retain_id_t0 = _1012_ | _1011_;
  assign perf_tbranch_o_t0 = _1015_ | _1014_;
  assign perf_jump_o_t0 = _1017_ | _1016_;
  assign debug_cause_o_t0 = _1021_ | _1434_;
  assign csr_mtval_o_t0 = _1024_ | _1437_;
  assign csr_restore_dret_id_o_t0 = _1026_ | _1025_;
  assign csr_restore_mret_id_o_t0 = _1028_ | _1027_;
  assign csr_save_wb_o_t0 = _1030_ | _1029_;
  assign _0019_ = _1038_ | _1440_;
  assign _0015_ = _1041_ | _1443_;
  assign _0011_ = _1044_ | _1446_;
  assign _0007_ = _1047_ | _1449_;
  assign _0003_ = _1050_ | _1452_;
  assign _0178_ = _1053_ | _1455_;
  assign _0172_ = _1056_ | _1458_;
  assign _0164_ = _1059_ | _1461_;
  assign _0156_ = _1062_ | _1464_;
  assign _0144_ = _1065_ | _1467_;
  assign _0126_ = _1068_ | _1470_;
  assign _0103_ = _1071_ | _1473_;
  assign _0062_ = _1074_ | _1476_;
  assign mfip_id_t0 = _1077_ | _1479_;
  assign do_single_step_d_t0 = _1080_ | _1482_;
  assign _1769_ = _1082_ | _1081_;
  assign ebreak_into_debug_t0 = _1085_ | _1486_;
  assign _1771_ = _1088_ | _1489_;
  assign _1773_ = _1091_ | _1492_;
  assign _1775_ = _1094_ | _1495_;
  assign _1777_ = _1097_ | _1498_;
  assign _0193_ = { _1719_, _1686_, dret_insn, mret_insn } != 4'h8;
  assign _0195_ = { _1719_, _1686_, mret_insn } != 3'h5;
  assign _0197_ = { _1719_, _1686_ } != 2'h3;
  assign _0199_ = | { _0219_, _1719_ };
  assign _0201_ = { _1719_, _1686_, mret_insn } != 3'h4;
  assign _0203_ = { _1759_, handle_irq } != 2'h2;
  assign _0205_ = { _1759_, _1657_, handle_irq } != 3'h5;
  assign _0207_ = | { _1719_, _1759_ };
  assign _0209_ = { _1761_, id_in_ready_o, handle_irq, enter_debug_mode } != 4'h8;
  assign _0211_ = { _1762_, _1677_ } != 2'h2;
  assign _0213_ = & { _0197_, _0199_, _0193_, _0195_ };
  assign _0215_ = & { _0207_, _0203_, _0197_, _0201_, _0205_ };
  assign _0217_ = & { _0209_, _0211_ };
  assign _0410_ = ~ _0034_;
  assign _0411_ = ~ _0122_;
  assign _0412_ = ~ _0161_;
  assign _0413_ = ~ _0141_;
  assign _0414_ = ~ _0045_;
  assign _0415_ = ~ _0107_;
  assign _0417_ = ~ _1744_;
  assign _0418_ = ~ _1746_;
  assign _0419_ = ~ _1748_;
  assign _0420_ = ~ _0130_;
  assign _0421_ = ~ _0095_;
  assign _0422_ = ~ _1639_;
  assign _0221_ = | { _1766_, _1764_, _1758_, _1756_ };
  assign _0223_ = | { _1763_, _1762_, _1758_, _1756_ };
  assign _0227_ = | { _1764_, _1761_, _1760_, _1759_, _1758_, _1756_, _1719_ };
  assign _0225_ = | { _1759_, _1758_, _1756_ };
  assign _0228_ = | { _1763_, _1762_, _1719_ };
  assign _0251_ = ~ _0221_;
  assign _0253_ = ~ _0225_;
  assign _0302_ = ~ illegal_insn_i;
  assign _0304_ = ~ _1697_;
  assign _0308_ = ~ _1701_;
  assign _0310_ = ~ _1703_;
  assign _0314_ = ~ wfi_insn;
  assign _0317_ = ~ _1707_;
  assign _0319_ = ~ _1709_;
  assign _0321_ = ~ special_req_pc_change;
  assign _0110_ = ~ _0082_;
  assign _0324_ = ~ _1711_;
  assign _0282_ = ~ debug_req_i;
  assign _0326_ = ~ enter_debug_mode_prio_d;
  assign _0279_ = ~ irq_nm_i;
  assign _0329_ = ~ ready_wb_i;
  assign _0284_ = ~ debug_mode_o;
  assign _0332_ = ~ stall_id_i;
  assign _0292_ = ~ stall;
  assign _0301_ = ~ _0181_;
  assign _0303_ = ~ illegal_dret;
  assign _0305_ = ~ illegal_umode;
  assign _0309_ = ~ illegal_insn_d;
  assign _0315_ = ~ csr_pipe_flush;
  assign _0318_ = ~ exc_req_d;
  assign _0320_ = ~ exc_req_lsu;
  assign _0322_ = ~ special_req_flush_only;
  assign _0313_ = ~ load_err_i;
  assign _0312_ = ~ store_err_i;
  assign _0325_ = ~ do_single_step_d;
  assign _0327_ = ~ _0185_;
  assign _0328_ = ~ _0189_;
  assign _0330_ = ~ wb_exception_o;
  assign _0331_ = ~ ebreak_into_debug;
  assign _0333_ = ~ stall_wb_i;
  assign _0334_ = ~ retain_id;
  assign _0336_ = ~ flush_id_o;
  assign _0555_ = _0659_ & _0250_;
  assign _0558_ = _0222_ & _0252_;
  assign _0561_ = _0226_ & _0252_;
  assign _0564_ = controller_run_o_t0 & _0255_;
  assign _0567_ = _1757_ & _0252_;
  assign _0722_ = mret_insn_t0 & _0301_;
  assign _0725_ = illegal_insn_i_t0 & _0303_;
  assign _0728_ = _1698_ & _0305_;
  assign _0731_ = ecall_insn_t0 & _0307_;
  assign _0734_ = _1702_ & _0309_;
  assign _0737_ = _1704_ & _0311_;
  assign _0740_ = store_err_i_t0 & _0313_;
  assign _0743_ = wfi_insn_t0 & _0315_;
  assign _0746_ = mret_insn_t0 & _0316_;
  assign _0749_ = _1708_ & _0318_;
  assign _0752_ = _1710_ & _0320_;
  assign _0755_ = special_req_pc_change_t0 & _0322_;
  assign _0758_ = instr_valid_i_t0 & ready_wb_i;
  assign _0761_ = load_err_q_t0 & _0295_;
  assign _0764_ = _0083_ & _0313_;
  assign _0767_ = _1712_ & _0312_;
  assign _0770_ = debug_req_i_t0 & _0325_;
  assign _0773_ = enter_debug_mode_prio_d_t0 & _0327_;
  assign _0776_ = irq_nm_i_t0 & _0328_;
  assign _0779_ = ready_wb_i_t0 & _0330_;
  assign _0782_ = debug_mode_o_t0 & _0331_;
  assign _0784_ = stall_id_i_t0 & _0333_;
  assign _0787_ = stall_t0 & _0334_;
  assign _0790_ = _1694_ & _0336_;
  assign _0556_ = _1145_[1] & _0249_;
  assign _0559_ = _1141_[3] & _0251_;
  assign _0562_ = _1141_[3] & _0253_;
  assign _0565_ = _0229_ & _0254_;
  assign _0568_ = _1141_[3] & _0256_;
  assign _0723_ = _0182_ & _0300_;
  assign _0726_ = illegal_dret_t0 & _0302_;
  assign _0729_ = illegal_umode_t0 & _0304_;
  assign _0732_ = ebrk_insn_t0 & _0306_;
  assign _0735_ = illegal_insn_d_t0 & _0308_;
  assign _0738_ = instr_fetch_err_t0 & _0310_;
  assign _0741_ = load_err_i_t0 & _0312_;
  assign _0744_ = csr_pipe_flush_t0 & _0314_;
  assign _0747_ = dret_insn_t0 & _0300_;
  assign _0750_ = exc_req_d_t0 & _0317_;
  assign _0753_ = exc_req_lsu_t0 & _0319_;
  assign _0756_ = special_req_flush_only_t0 & _0321_;
  assign _0759_ = ready_wb_i_t0 & _0323_;
  assign _0762_ = store_err_prio_t0 & _0297_;
  assign _0765_ = load_err_i_t0 & _0110_;
  assign _0768_ = store_err_i_t0 & _0324_;
  assign _0771_ = do_single_step_d_t0 & _0282_;
  assign _0774_ = _0186_ & _0326_;
  assign _0777_ = _0190_ & _0279_;
  assign _0780_ = wb_exception_o_t0 & _0329_;
  assign _0783_ = ebreak_into_debug_t0 & _0284_;
  assign _0785_ = stall_wb_i_t0 & _0332_;
  assign _0788_ = retain_id_t0 & _0292_;
  assign _0791_ = flush_id_o_t0 & _0335_;
  assign _0557_ = _0659_ & _1145_[1];
  assign _0560_ = _0222_ & _1141_[3];
  assign _0563_ = _0226_ & _1141_[3];
  assign _0566_ = controller_run_o_t0 & _0229_;
  assign _0569_ = _1757_ & _1141_[3];
  assign _0724_ = mret_insn_t0 & _0182_;
  assign _0727_ = illegal_insn_i_t0 & illegal_dret_t0;
  assign _0730_ = _1698_ & illegal_umode_t0;
  assign _0733_ = ecall_insn_t0 & ebrk_insn_t0;
  assign _0736_ = _1702_ & illegal_insn_d_t0;
  assign _0739_ = _1704_ & instr_fetch_err_t0;
  assign _0742_ = store_err_i_t0 & load_err_i_t0;
  assign _0745_ = wfi_insn_t0 & csr_pipe_flush_t0;
  assign _0748_ = mret_insn_t0 & dret_insn_t0;
  assign _0751_ = _1708_ & exc_req_d_t0;
  assign _0754_ = _1710_ & exc_req_lsu_t0;
  assign _0757_ = special_req_pc_change_t0 & special_req_flush_only_t0;
  assign _0760_ = instr_valid_i_t0 & ready_wb_i_t0;
  assign _0763_ = load_err_q_t0 & store_err_prio_t0;
  assign _0766_ = _0083_ & load_err_i_t0;
  assign _0769_ = _1712_ & store_err_i_t0;
  assign _0772_ = debug_req_i_t0 & do_single_step_d_t0;
  assign _0775_ = enter_debug_mode_prio_d_t0 & _0186_;
  assign _0778_ = irq_nm_i_t0 & _0190_;
  assign _0781_ = ready_wb_i_t0 & wb_exception_o_t0;
  assign _0679_ = debug_mode_o_t0 & ebreak_into_debug_t0;
  assign _0786_ = stall_id_i_t0 & stall_wb_i_t0;
  assign _0789_ = stall_t0 & retain_id_t0;
  assign _0792_ = _1694_ & flush_id_o_t0;
  assign _1149_ = _0555_ | _0556_;
  assign _1150_ = _0558_ | _0559_;
  assign _1151_ = _0561_ | _0562_;
  assign _1152_ = _0564_ | _0565_;
  assign _1153_ = _0567_ | _0568_;
  assign _1246_ = _0722_ | _0723_;
  assign _1247_ = _0725_ | _0726_;
  assign _1248_ = _0728_ | _0729_;
  assign _1249_ = _0731_ | _0732_;
  assign _1250_ = _0734_ | _0735_;
  assign _1251_ = _0737_ | _0738_;
  assign _1252_ = _0740_ | _0741_;
  assign _1253_ = _0743_ | _0744_;
  assign _1254_ = _0746_ | _0747_;
  assign _1255_ = _0749_ | _0750_;
  assign _1256_ = _0752_ | _0753_;
  assign _1257_ = _0755_ | _0756_;
  assign _1258_ = _0758_ | _0759_;
  assign _1259_ = _0761_ | _0762_;
  assign _1260_ = _0764_ | _0765_;
  assign _1261_ = _0767_ | _0768_;
  assign _1262_ = _0770_ | _0771_;
  assign _1263_ = _0773_ | _0774_;
  assign _1264_ = _0776_ | _0777_;
  assign _1265_ = _0779_ | _0780_;
  assign _1266_ = _0782_ | _0783_;
  assign _1267_ = _0784_ | _0785_;
  assign _1268_ = _0787_ | _0788_;
  assign _1269_ = _0790_ | _0791_;
  assign _1101_ = _1149_ | _0557_;
  assign _1103_ = _1150_ | _0560_;
  assign _1099_ = _1151_ | _0563_;
  assign _1105_ = _1152_ | _0566_;
  assign _1107_ = _1153_ | _0569_;
  assign _1696_ = _1246_ | _0724_;
  assign _1698_ = _1247_ | _0727_;
  assign _1700_ = _1248_ | _0730_;
  assign _1702_ = _1249_ | _0733_;
  assign _1704_ = _1250_ | _0736_;
  assign _1706_ = _1251_ | _0739_;
  assign exc_req_lsu_t0 = _1252_ | _0742_;
  assign special_req_flush_only_t0 = _1253_ | _0745_;
  assign _1708_ = _1254_ | _0748_;
  assign _1710_ = _1255_ | _0751_;
  assign special_req_pc_change_t0 = _1256_ | _0754_;
  assign special_req_t0 = _1257_ | _0757_;
  assign id_wb_pending_t0 = _1258_ | _0760_;
  assign _0083_ = _1259_ | _0763_;
  assign _1712_ = _1260_ | _0766_;
  assign wb_exception_o_t0 = _1261_ | _0769_;
  assign _1714_ = _1262_ | _0772_;
  assign enter_debug_mode_t0 = _1263_ | _0775_;
  assign _1716_ = _1264_ | _0778_;
  assign _1718_ = _1265_ | _0781_;
  assign _0121_ = _1266_ | _0679_;
  assign stall_t0 = _1267_ | _0786_;
  assign _1694_ = _1268_ | _0789_;
  assign instr_valid_clear_o_t0 = _1269_ | _0792_;
  assign _0219_ = | { _1758_, _1756_ };
  assign _1100_ = _1763_ | _1762_;
  assign _1102_ = _0221_ | _1719_;
  assign _1098_ = _0225_ | _1719_;
  assign _1104_ = _1760_ | _0228_;
  assign _1106_ = _1756_ | _1719_;
  assign _0426_ = | { _1761_, _1760_, _1098_ };
  assign _1603_ = _1719_ ? _0026_ : 4'h5;
  assign _1605_ = _1760_ ? _0167_ : _0134_;
  assign _1607_ = _1098_ ? _1603_ : _1605_;
  assign _1609_ = _1762_ ? _0041_ : 4'h3;
  assign _1611_ = _1766_ ? 4'h1 : 4'h0;
  assign _1613_ = _1764_ ? 4'h4 : _1611_;
  assign _1615_ = _1100_ ? _1609_ : _1613_;
  assign ctrl_fsm_ns = _0426_ ? _1607_ : _1615_;
  assign _1619_ = _1760_ ? _0068_ : 1'h0;
  assign _1621_ = _1759_ ? _0034_ : _1619_;
  assign pc_set_spec_o = _1102_ ? _1617_ : _1621_;
  assign _1617_ = _1719_ ? _0130_ : 1'h1;
  assign _1623_ = _1760_ ? _0066_ : 1'h0;
  assign _1625_ = _1759_ ? _0034_ : _1623_;
  assign pc_set_o = _1102_ ? _1617_ : _1625_;
  assign _1627_ = _1719_ ? _0064_ : 3'h2;
  assign _1629_ = _1760_ ? 3'h1 : 3'h0;
  assign pc_mux_o = _1098_ ? _1627_ : _1629_;
  assign _1631_ = _0228_ ? 1'h1 : _0141_;
  assign _1633_ = _1761_ ? _0097_ : 1'h0;
  assign halt_if = _1104_ ? _1631_ : _1633_;
  assign debug_mode_d = _1719_ ? _0045_ : 1'h1;
  assign nmi_mode_d = _1719_ ? _0127_ : _0063_;
  assign _1635_ = _0223_ ? 1'h1 : 1'h0;
  assign flush_id_o = _1719_ ? _0054_ : _1635_;
  assign _1636_ = _1758_ ? 1'h1 : 1'h0;
  assign debug_csr_save_o = _1756_ ? _0035_ : _1636_;
  assign _1637_ = _1719_ ? _0108_ : _0035_;
  assign csr_save_if_o = _1758_ ? 1'h1 : _1639_;
  assign csr_save_cause_o = _1106_ ? _1637_ : csr_save_if_o;
  assign _1641_ = _1756_ ? _0035_ : 1'h0;
  assign csr_save_id_o = _1719_ ? _0080_ : _1641_;
  assign _1639_ = _1759_ ? _0034_ : 1'h0;
  assign _1643_ = _1759_ ? _0050_ : 6'h00;
  assign exc_cause_o = _1719_ ? _0159_ : _1643_;
  assign _1645_ = _0219_ ? 2'h2 : 2'h1;
  assign exc_pc_mux_o = _1719_ ? _0052_ : _1645_;
  assign _1647_ = _1763_ ? 1'h0 : 1'h1;
  assign ctrl_busy_o = _1762_ ? _0039_ : _1647_;
  assign _0437_ = | { _0200_, _0198_, _0196_, _0194_ };
  assign _0438_ = | { _0208_, _0206_, _0204_, _0202_, _0198_ };
  assign _0439_ = | { _0212_, _0210_ };
  assign _1146_ = { _0197_, _0199_, _0193_, _0195_ } | { _0198_, _0200_, _0194_, _0196_ };
  assign _1147_ = { _0207_, _0203_, _0197_, _0201_, _0205_ } | { _0208_, _0204_, _0198_, _0202_, _0206_ };
  assign _1148_ = { _0209_, _0211_ } | { _0210_, _0212_ };
  assign _0423_ = & _1146_;
  assign _0424_ = & _1147_;
  assign _0425_ = & _1148_;
  assign _0214_ = _0437_ & _0423_;
  assign _0216_ = _0438_ & _0424_;
  assign _0218_ = _0439_ & _0425_;
  assign _1650_ = ! priv_mode_i;
  assign _1648_ = priv_mode_i == 2'h3;
  assign _1652_ = _1680_ && _1682_;
  assign _1653_ = _1665_ && _1666_;
  assign _1655_ = _1653_ && _1667_;
  assign _1657_ = irq_nm_i && _1668_;
  assign _1658_ = ebreak_into_debug && _1669_;
  assign _1659_ = csr_pipe_flush && handle_irq;
  assign _1661_ = ebrk_insn_prio && ebreak_into_debug;
  assign _1663_ = enter_debug_mode_prio_q && _1670_;
  assign _1665_ = ! stall;
  assign _1666_ = ! special_req;
  assign _1667_ = ! id_wb_pending;
  assign _1668_ = ! nmi_mode_o;
  assign _1669_ = ! debug_mode_o;
  assign _1670_ = ! _1661_;
  assign _1671_ = irq_nm_i || irq_pending_i;
  assign _1673_ = _1671_ || debug_req_i;
  assign _1675_ = _1673_ || debug_mode_o;
  assign _1677_ = _1675_ || debug_single_step_i;
  assign _1678_ = branch_set_i || jump_set_i;
  assign _1679_ = branch_set_spec_i || jump_set_i;
  assign _1680_ = enter_debug_mode || handle_irq;
  assign _1682_ = stall || id_wb_pending;
  assign _1684_ = exc_req_q || store_err_q;
  assign _1686_ = _1684_ || load_err_q;
  assign _1687_ = priv_mode_i != 2'h3;
  assign _1688_ = ctrl_fsm_cs != 4'h6;
  assign _1689_ = | irqs_i[14:0];
  assign _1691_ = ~ nmi_mode_o;
  assign _1692_ = ~ halt_if;
  assign _1693_ = ~ _0335_;
  assign _1695_ = mret_insn | _0181_;
  assign _1697_ = illegal_insn_i | illegal_dret;
  assign _1699_ = _1697_ | illegal_umode;
  assign _1701_ = ecall_insn | ebrk_insn;
  assign _1703_ = _1701_ | illegal_insn_d;
  assign _1705_ = _1703_ | instr_fetch_err;
  assign exc_req_lsu = store_err_i | load_err_i;
  assign special_req_flush_only = wfi_insn | csr_pipe_flush;
  assign _1707_ = mret_insn | dret_insn;
  assign _1709_ = _1707_ | exc_req_d;
  assign special_req_pc_change = _1709_ | exc_req_lsu;
  assign special_req = special_req_pc_change | special_req_flush_only;
  assign id_wb_pending = instr_valid_i | _0329_;
  assign _0082_ = load_err_q | store_err_q;
  assign _1711_ = _0082_ | load_err_i;
  assign wb_exception_o = _1711_ | store_err_i;
  assign _1713_ = debug_req_i | do_single_step_d;
  assign enter_debug_mode = enter_debug_mode_prio_d | _0185_;
  assign _1715_ = irq_nm_i | _0189_;
  assign _1717_ = ready_wb_i | wb_exception_o;
  assign _0416_ = debug_mode_o | ebreak_into_debug;
  assign stall = stall_id_i | stall_wb_i;
  assign _0335_ = stall | retain_id;
  assign instr_valid_clear_o = _1693_ | flush_id_o;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) load_err_q <= 1'h0;
    else load_err_q <= load_err_i;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) store_err_q <= 1'h0;
    else store_err_q <= store_err_i;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) exc_req_q <= 1'h0;
    else exc_req_q <= exc_req_d;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) illegal_insn_q <= 1'h0;
    else illegal_insn_q <= illegal_insn_d;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) do_single_step_q <= 1'h0;
    else do_single_step_q <= do_single_step_d;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) enter_debug_mode_prio_q <= 1'h0;
    else enter_debug_mode_prio_q <= enter_debug_mode_prio_d;
  assign _0150_ = ebrk_insn ? 1'h1 : 1'h0;
  assign _0138_ = ecall_insn ? 1'h1 : 1'h0;
  assign _0136_ = ecall_insn ? 1'h0 : _0150_;
  assign _0124_ = illegal_insn_q ? 1'h1 : 1'h0;
  assign _0114_ = illegal_insn_q ? 1'h0 : _0136_;
  assign _0116_ = illegal_insn_q ? 1'h0 : _0138_;
  assign _0101_ = instr_fetch_err ? 1'h1 : 1'h0;
  assign _0089_ = instr_fetch_err ? 1'h0 : _0114_;
  assign _0091_ = instr_fetch_err ? 1'h0 : _0116_;
  assign _0099_ = instr_fetch_err ? 1'h0 : _0124_;
  assign _0060_ = load_err_q ? 1'h1 : 1'h0;
  assign _0046_ = load_err_q ? 1'h0 : _0089_;
  assign _0048_ = load_err_q ? 1'h0 : _0091_;
  assign _0056_ = load_err_q ? 1'h0 : _0099_;
  assign _0058_ = load_err_q ? 1'h0 : _0101_;
  assign store_err_prio = store_err_q ? 1'h1 : 1'h0;
  assign load_err_prio = store_err_q ? 1'h0 : _0060_;
  assign ebrk_insn_prio = store_err_q ? 1'h0 : _0046_;
  assign ecall_insn_prio = store_err_q ? 1'h0 : _0048_;
  assign illegal_insn_prio = store_err_q ? 1'h0 : _0056_;
  assign instr_fetch_err_prio = store_err_q ? 1'h0 : _0058_;
  assign _0026_ = _1663_ ? 4'h8 : _0004_;
  assign _0024_ = _1659_ ? 4'h7 : 4'h5;
  assign _0022_ = wfi_insn ? 4'h2 : _0024_;
  assign _0113_ = dret_insn ? 1'h0 : 1'hx;
  assign _0107_ = dret_insn ? 1'h1 : 1'h0;
  assign _0128_ = dret_insn ? 3'h4 : 3'h0;
  assign _0020_ = dret_insn ? 4'h5 : _0022_;
  assign _0145_ = mret_insn ? 1'h0 : 1'hx;
  assign _0079_ = mret_insn ? 1'h1 : 1'h0;
  assign _0165_ = mret_insn ? 1'h1 : _0107_;
  assign _0105_ = mret_insn ? 3'h3 : _0128_;
  assign _0088_ = mret_insn ? 1'hx : _0113_;
  assign _0016_ = mret_insn ? 4'h5 : _0020_;
  assign _0077_ = mret_insn ? 1'h0 : _0107_;
  assign _0012_ = _0416_ ? 4'h9 : 4'h5;
  assign _0120_ = _0416_ ? 1'h0 : 1'h1;
  assign _0146_ = _0416_ ? 1'h0 : _0110_;
  assign _0175_ = _0416_ ? 6'h00 : 6'h03;
  assign _1720_ = load_err_prio ? lsu_addr_last_i : 32'd0;
  assign _1532_ = store_err_prio ? lsu_addr_last_i : _1720_;
  assign _1533_ = ebrk_insn_prio ? 32'd0 : _1532_;
  assign _1724_ = ecall_insn_prio ? 32'd0 : _1533_;
  assign _1726_ = illegal_insn_prio ? _1774_ : _1724_;
  assign _0075_ = instr_fetch_err_prio ? _1772_ : _1726_;
  assign _1728_ = load_err_prio ? 6'h05 : 6'h00;
  assign _1730_ = store_err_prio ? 6'h07 : _1728_;
  assign _1732_ = ebrk_insn_prio ? _0175_ : _1730_;
  assign _1734_ = ecall_insn_prio ? _1776_ : _1732_;
  assign _1736_ = illegal_insn_prio ? 6'h02 : _1734_;
  assign _0169_ = instr_fetch_err_prio ? 6'h01 : _1736_;
  assign _1738_ = ebrk_insn_prio ? _0012_ : 4'h5;
  assign _1740_ = ecall_insn_prio ? 4'h5 : _1738_;
  assign _1742_ = illegal_insn_prio ? 4'h5 : _1740_;
  assign _0008_ = instr_fetch_err_prio ? 4'h5 : _1742_;
  assign _1748_ = illegal_insn_prio ? 1'h1 : _1746_;
  assign _0095_ = instr_fetch_err_prio ? 1'h1 : _1748_;
  assign _1750_ = ebrk_insn_prio ? _0146_ : _0110_;
  assign _1752_ = ecall_insn_prio ? _0110_ : _1750_;
  assign _1754_ = illegal_insn_prio ? _0110_ : _1752_;
  assign _0132_ = instr_fetch_err_prio ? _0110_ : _1754_;
  assign _1744_ = ebrk_insn_prio ? _0120_ : 1'h1;
  assign _1746_ = ecall_insn_prio ? 1'h1 : _1744_;
  assign _0004_ = _1686_ ? _0008_ : _0016_;
  assign _0054_ = _1686_ ? _0095_ : 1'h1;
  assign _0028_ = _1686_ ? _0075_ : 32'd0;
  assign _0108_ = _1686_ ? _0095_ : 1'h0;
  assign _0080_ = _1686_ ? _0132_ : 1'h0;
  assign _0159_ = _1686_ ? _0169_ : 6'h00;
  assign _0130_ = _1686_ ? _0095_ : _0165_;
  assign _0037_ = _1686_ ? _0082_ : 1'h0;
  assign _0052_ = _1686_ ? _1770_ : 2'h1;
  assign _0064_ = _1686_ ? 3'h2 : _0105_;
  assign _0045_ = _1686_ ? 1'hx : _0088_;
  assign _0127_ = _1686_ ? 1'hx : _0145_;
  assign _0030_ = _1686_ ? 1'h0 : _0077_;
  assign _0032_ = _1686_ ? 1'h0 : _0079_;
  assign _0035_ = _1658_ ? 1'h1 : 1'h0;
  assign _0086_ = debug_single_step_i ? 3'h4 : 3'h3;
  assign _0043_ = trigger_match_i ? 3'h2 : _0086_;
  assign _0151_ = irqs_i[17] ? 6'h23 : 6'h27;
  assign _0139_ = irqs_i[15] ? 6'h2b : _0151_;
  assign _0118_ = _1689_ ? { 2'h3, mfip_id } : _0139_;
  assign _0104_ = _1657_ ? 1'h1 : 1'hx;
  assign _0093_ = _1657_ ? 6'h3f : _0118_;
  assign _0063_ = handle_irq ? _0104_ : 1'hx;
  assign _0050_ = handle_irq ? _0093_ : 6'h00;
  assign _0034_ = handle_irq ? 1'h1 : 1'h0;
  assign _0161_ = handle_irq ? 1'h1 : _0122_;
  assign _0000_ = handle_irq ? 4'h7 : _0148_;
  assign _0153_ = enter_debug_mode ? 1'h1 : _0161_;
  assign _0173_ = enter_debug_mode ? 4'h8 : _0000_;
  assign _0141_ = _1655_ ? _0153_ : _0122_;
  assign _0167_ = _1655_ ? _0173_ : _0148_;
  assign _0122_ = _1652_ ? 1'h1 : 1'h0;
  assign _0068_ = _1679_ ? 1'h1 : 1'h0;
  assign _0070_ = _1678_ ? jump_set_i : 1'h0;
  assign _0072_ = _1678_ ? branch_set_i : 1'h0;
  assign _0066_ = _1678_ ? 1'h1 : 1'h0;
  assign _0157_ = _1717_ ? 4'h6 : ctrl_fsm_cs;
  assign _0148_ = special_req ? _0157_ : ctrl_fsm_cs;
  assign _0074_ = special_req ? 1'h1 : 1'h0;
  assign _0097_ = enter_debug_mode ? 1'h1 : _0034_;
  assign _0134_ = enter_debug_mode ? 4'h8 : _0111_;
  assign _0111_ = handle_irq ? 4'h7 : _0084_;
  assign _0084_ = id_in_ready_o ? 4'h5 : 4'hx;
  assign _0041_ = _1677_ ? 4'h4 : 4'hx;
  assign _0039_ = _1677_ ? 1'h1 : 1'h0;
  assign _1766_ = ! ctrl_fsm_cs;
  assign instr_req_o = _0227_ ? 1'h1 : 1'h0;
  assign _1764_ = ctrl_fsm_cs == 4'h1;
  assign retain_id = _1760_ ? _0074_ : 1'h0;
  assign _1761_ = ctrl_fsm_cs == 4'h4;
  assign controller_run_o = _1760_ ? 1'h1 : 1'h0;
  assign perf_tbranch_o = _1760_ ? _0072_ : 1'h0;
  assign perf_jump_o = _1760_ ? _0070_ : 1'h0;
  assign _1760_ = ctrl_fsm_cs == 4'h5;
  assign debug_cause_o = _1758_ ? _0043_ : 3'h1;
  assign csr_mtval_o = _1719_ ? _0028_ : 32'd0;
  assign csr_restore_dret_id_o = _1719_ ? _0030_ : 1'h0;
  assign csr_restore_mret_id_o = _1719_ ? _0032_ : 1'h0;
  assign csr_save_wb_o = _1719_ ? _0037_ : 1'h0;
  assign _1759_ = ctrl_fsm_cs == 4'h7;
  assign _1719_ = ctrl_fsm_cs == 4'h6;
  assign _1756_ = ctrl_fsm_cs == 4'h9;
  assign _1758_ = ctrl_fsm_cs == 4'h8;
  assign _1762_ = ctrl_fsm_cs == 4'h3;
  assign _1763_ = ctrl_fsm_cs == 4'h2;
  assign _0018_ = irqs_i[1] ? 4'h1 : 4'h0;
  assign _0014_ = irqs_i[2] ? 4'h2 : _0018_;
  assign _0010_ = irqs_i[3] ? 4'h3 : _0014_;
  assign _0006_ = irqs_i[4] ? 4'h4 : _0010_;
  assign _0002_ = irqs_i[5] ? 4'h5 : _0006_;
  assign _0177_ = irqs_i[6] ? 4'h6 : _0002_;
  assign _0171_ = irqs_i[7] ? 4'h7 : _0177_;
  assign _0163_ = irqs_i[8] ? 4'h8 : _0171_;
  assign _0155_ = irqs_i[9] ? 4'h9 : _0163_;
  assign _0143_ = irqs_i[10] ? 4'ha : _0155_;
  assign _0125_ = irqs_i[11] ? 4'hb : _0143_;
  assign _0102_ = irqs_i[12] ? 4'hc : _0125_;
  assign _0061_ = irqs_i[13] ? 4'hd : _0102_;
  assign mfip_id = irqs_i[14] ? 4'he : _0061_;
  assign do_single_step_d = instr_valid_i ? _0183_ : do_single_step_q;
  assign _1768_ = _1650_ ? debug_ebreaku_i : 1'h0;
  assign ebreak_into_debug = _1648_ ? debug_ebreakm_i : _1768_;
  assign _1770_ = debug_mode_o ? 2'h3 : 2'h0;
  assign _1772_ = instr_fetch_err_plus2_i ? _0179_ : pc_id_i;
  assign _1774_ = instr_is_compressed_i ? { 16'h0000, instr_compressed_i } : instr_i;
  assign _1776_ = _1648_ ? 6'h0b : 6'h08;
  assign _1141_[1:0] = { dret_insn_t0, mret_insn_t0 };
  assign _1142_[0] = handle_irq_t0;
  assign { _1143_[2], _1143_[0] } = { _1142_[1], handle_irq_t0 };
  assign _1144_[2:0] = { id_in_ready_o_t0, handle_irq_t0, enter_debug_mode_t0 };
  assign _1145_[0] = _0040_;
  assign nt_branch_mispredict_o = 1'h0;
  assign nt_branch_mispredict_o_t0 = 1'h0;
endmodule

module paramodauxy_ibex_counterCounterWidth3200000000000000000000000000100000 (clk_i, rst_ni, counter_inc_i, counterh_we_i, counter_we_i, counter_val_i, counter_val_o, counter_inc_i_t0, counter_val_i_t0, counter_val_o_t0, counter_we_i_t0, counterh_we_i_t0);
  wire [31:0] _000_;
  wire [31:0] _001_;
  wire _002_;
  wire _003_;
  wire _004_;
  wire _005_;
  wire _006_;
  wire _007_;
  wire [31:0] _008_;
  wire _009_;
  wire [1:0] _010_;
  wire [1:0] _011_;
  wire _012_;
  wire _013_;
  wire [31:0] _014_;
  wire [31:0] _015_;
  wire [31:0] _016_;
  wire _017_;
  wire _018_;
  wire _019_;
  wire _020_;
  wire _021_;
  wire [31:0] _022_;
  wire [31:0] _023_;
  wire [31:0] _024_;
  wire [31:0] _025_;
  wire [1:0] _026_;
  wire [1:0] _027_;
  wire [1:0] _028_;
  wire _029_;
  wire _030_;
  wire _031_;
  wire [31:0] _032_;
  wire [31:0] _033_;
  wire [31:0] _034_;
  wire [31:0] _035_;
  wire [31:0] _036_;
  wire [31:0] _037_;
  wire [31:0] _038_;
  wire [31:0] _039_;
  wire [31:0] _040_;
  wire [31:0] _041_;
  wire [31:0] _042_;
  wire [31:0] _043_;
  wire [31:0] _044_;
  wire [31:0] _045_;
  wire [1:0] _046_;
  wire _047_;
  wire [31:0] _048_;
  wire [31:0] _049_;
  wire [31:0] _050_;
  wire [31:0] _051_;
  wire [31:0] _052_;
  wire [31:0] _053_;
  wire [31:0] _054_;
  wire [31:0] _055_;
  wire [31:0] _056_;
  wire [31:0] _057_;
  wire [31:0] _058_;
  wire [31:0] _059_;
  wire _060_;
  wire [31:0] _061_;
  wire [31:0] _062_;
  input clk_i;
  wire clk_i;
  wire [31:0] counter_d;
  wire [31:0] counter_d_t0;
  input counter_inc_i;
  wire counter_inc_i;
  input counter_inc_i_t0;
  wire counter_inc_i_t0;
  wire [63:0] counter_load;
  wire [63:0] counter_load_t0;
  reg [31:0] counter_q;
  reg [31:0] counter_q_t0;
  wire [31:0] counter_upd;
  wire [31:0] counter_upd_t0;
  input [31:0] counter_val_i;
  wire [31:0] counter_val_i;
  input [31:0] counter_val_i_t0;
  wire [31:0] counter_val_i_t0;
  output [63:0] counter_val_o;
  wire [63:0] counter_val_o;
  output [63:0] counter_val_o_t0;
  wire [63:0] counter_val_o_t0;
  input counter_we_i;
  wire counter_we_i;
  input counter_we_i_t0;
  wire counter_we_i_t0;
  input counterh_we_i;
  wire counterh_we_i;
  input counterh_we_i_t0;
  wire counterh_we_i_t0;
  input rst_ni;
  wire rst_ni;
  wire we;
  wire we_t0;
  assign counter_upd = counter_q + 32'd1;
  assign _008_ = ~ counter_q_t0;
  assign _022_ = counter_q & _008_;
  assign _061_ = _022_ + 32'd1;
  assign _041_ = counter_q | counter_q_t0;
  assign _062_ = _041_ + 32'd1;
  assign _057_ = _061_ ^ _062_;
  assign counter_upd_t0 = _057_ | counter_q_t0;
  assign _009_ = ~ _006_;
  assign _058_ = counter_d ^ counter_q;
  assign _042_ = counter_d_t0 | counter_q_t0;
  assign _043_ = _058_ | _042_;
  assign _023_ = { _006_, _006_, _006_, _006_, _006_, _006_, _006_, _006_, _006_, _006_, _006_, _006_, _006_, _006_, _006_, _006_, _006_, _006_, _006_, _006_, _006_, _006_, _006_, _006_, _006_, _006_, _006_, _006_, _006_, _006_, _006_, _006_ } & counter_d_t0;
  assign _024_ = { _009_, _009_, _009_, _009_, _009_, _009_, _009_, _009_, _009_, _009_, _009_, _009_, _009_, _009_, _009_, _009_, _009_, _009_, _009_, _009_, _009_, _009_, _009_, _009_, _009_, _009_, _009_, _009_, _009_, _009_, _009_, _009_ } & counter_q_t0;
  assign _025_ = _043_ & { _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_ };
  assign _044_ = _023_ | _024_;
  assign _045_ = _044_ | _025_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) counter_q_t0 <= 32'd0;
    else counter_q_t0 <= _045_;
  assign _019_ = | { we_t0, counterh_we_i_t0 };
  assign _011_ = ~ { we_t0, counterh_we_i_t0 };
  assign _027_ = { we, counterh_we_i } & _011_;
  assign _028_ = 2'h3 & _011_;
  assign _060_ = _027_ == _028_;
  assign _005_ = _060_ & _019_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) counter_q <= 32'd0;
    else if (_006_) counter_q <= counter_d;
  assign _018_ = | { we_t0, counter_inc_i_t0 };
  assign _010_ = ~ { we_t0, counter_inc_i_t0 };
  assign _026_ = { we, counter_inc_i } & _010_;
  assign _021_ = ! _026_;
  assign _003_ = _021_ & _018_;
  assign _014_ = ~ { counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i };
  assign _015_ = ~ { we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we };
  assign _016_ = ~ { counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i };
  assign _048_ = { counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0 } | _014_;
  assign _051_ = { we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0 } | _015_;
  assign _054_ = { counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0 } | _016_;
  assign _049_ = { counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0 } | { counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i };
  assign _052_ = { we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0 } | { we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we };
  assign _055_ = { counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0 } | { counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i };
  assign _032_ = 32'd0 & _048_;
  assign _035_ = _001_ & _051_;
  assign _038_ = counter_val_i_t0 & _054_;
  assign _033_ = counter_upd_t0 & _049_;
  assign _036_ = counter_load_t0[31:0] & _052_;
  assign _039_ = 32'd0 & _055_;
  assign _050_ = _032_ | _033_;
  assign _053_ = _035_ | _036_;
  assign _056_ = _038_ | _039_;
  assign _059_ = _000_ ^ counter_load[31:0];
  assign _034_ = { counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0 } & counter_upd;
  assign _037_ = { we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0 } & _059_;
  assign _040_ = { counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0 } & counter_val_i;
  assign _001_ = _034_ | _050_;
  assign counter_d_t0 = _037_ | _053_;
  assign counter_load_t0[31:0] = _040_ | _056_;
  assign _002_ = | { we, counter_inc_i };
  assign _004_ = { we, counterh_we_i } != 2'h3;
  assign _006_ = & { _004_, _002_ };
  assign _012_ = ~ counter_we_i;
  assign _013_ = ~ counterh_we_i;
  assign _029_ = counter_we_i_t0 & _013_;
  assign _030_ = counterh_we_i_t0 & _012_;
  assign _031_ = counter_we_i_t0 & counterh_we_i_t0;
  assign _047_ = _029_ | _030_;
  assign we_t0 = _047_ | _031_;
  assign _020_ = | { _005_, _003_ };
  assign _046_ = { _004_, _002_ } | { _005_, _003_ };
  assign _017_ = & _046_;
  assign _007_ = _020_ & _017_;
  assign we = counter_we_i | counterh_we_i;
  assign _000_ = counter_inc_i ? counter_upd : 32'hxxxxxxxx;
  assign counter_d = we ? counter_load[31:0] : _000_;
  assign counter_load[31:0] = counterh_we_i ? 32'hxxxxxxxx : counter_val_i;
  assign counter_val_o = { 32'h00000000, counter_q };
  assign counter_val_o_t0 = { 32'h00000000, counter_q_t0 };
endmodule

module paramodauxy_ibex_counterCounterWidths3200000000000000000000000001000000 (clk_i, rst_ni, counter_inc_i, counterh_we_i, counter_we_i, counter_val_i, counter_val_o, counter_inc_i_t0, counter_val_i_t0, counter_val_o_t0, counter_we_i_t0, counterh_we_i_t0);
  wire [63:0] _000_;
  wire [63:0] _001_;
  wire _002_;
  wire _003_;
  wire _004_;
  wire _005_;
  wire _006_;
  wire _007_;
  wire _008_;
  wire _009_;
  wire _010_;
  wire _011_;
  wire [63:0] _012_;
  wire _013_;
  wire _014_;
  wire [1:0] _015_;
  wire [1:0] _016_;
  wire _017_;
  wire _018_;
  wire [63:0] _019_;
  wire [63:0] _020_;
  wire [31:0] _021_;
  wire _022_;
  wire _023_;
  wire _024_;
  wire _025_;
  wire _026_;
  wire _027_;
  wire _028_;
  wire [63:0] _029_;
  wire [31:0] _030_;
  wire [31:0] _031_;
  wire [31:0] _032_;
  wire [31:0] _033_;
  wire [31:0] _034_;
  wire [31:0] _035_;
  wire [1:0] _036_;
  wire [1:0] _037_;
  wire [1:0] _038_;
  wire [1:0] _039_;
  wire _040_;
  wire _041_;
  wire _042_;
  wire [63:0] _043_;
  wire [63:0] _044_;
  wire [63:0] _045_;
  wire [63:0] _046_;
  wire [63:0] _047_;
  wire [63:0] _048_;
  wire [31:0] _049_;
  wire [31:0] _050_;
  wire [31:0] _051_;
  wire [31:0] _052_;
  wire [31:0] _053_;
  wire [63:0] _054_;
  wire [31:0] _055_;
  wire [31:0] _056_;
  wire [31:0] _057_;
  wire [31:0] _058_;
  wire [31:0] _059_;
  wire [31:0] _060_;
  wire [31:0] _061_;
  wire [31:0] _062_;
  wire [1:0] _063_;
  wire [1:0] _064_;
  wire _065_;
  wire [63:0] _066_;
  wire [63:0] _067_;
  wire [63:0] _068_;
  wire [63:0] _069_;
  wire [63:0] _070_;
  wire [63:0] _071_;
  wire [31:0] _072_;
  wire [31:0] _073_;
  wire [31:0] _074_;
  wire [31:0] _075_;
  wire [63:0] _076_;
  wire [31:0] _077_;
  wire [31:0] _078_;
  wire [63:0] _079_;
  wire _080_;
  wire _081_;
  wire [63:0] _082_;
  wire [63:0] _083_;
  input clk_i;
  wire clk_i;
  wire [63:0] counter_d;
  wire [63:0] counter_d_t0;
  input counter_inc_i;
  wire counter_inc_i;
  input counter_inc_i_t0;
  wire counter_inc_i_t0;
  wire [63:0] counter_load;
  wire [63:0] counter_load_t0;
  wire [63:0] counter_upd;
  wire [63:0] counter_upd_t0;
  input [31:0] counter_val_i;
  wire [31:0] counter_val_i;
  input [31:0] counter_val_i_t0;
  wire [31:0] counter_val_i_t0;
  output [63:0] counter_val_o;
  reg [63:0] counter_val_o;
  output [63:0] counter_val_o_t0;
  reg [63:0] counter_val_o_t0;
  input counter_we_i;
  wire counter_we_i;
  input counter_we_i_t0;
  wire counter_we_i_t0;
  input counterh_we_i;
  wire counterh_we_i;
  input counterh_we_i_t0;
  wire counterh_we_i_t0;
  input rst_ni;
  wire rst_ni;
  wire we;
  wire we_t0;
  assign counter_upd = counter_val_o + 64'h0000000000000001;
  assign _012_ = ~ counter_val_o_t0;
  assign _029_ = counter_val_o & _012_;
  assign _082_ = _029_ + 64'h0000000000000001;
  assign _054_ = counter_val_o | counter_val_o_t0;
  assign _083_ = _054_ + 64'h0000000000000001;
  assign _076_ = _082_ ^ _083_;
  assign counter_upd_t0 = _076_ | counter_val_o_t0;
  assign _013_ = ~ _008_;
  assign _014_ = ~ _010_;
  assign _077_ = counter_d[63:32] ^ counter_val_o[63:32];
  assign _078_ = counter_d[31:0] ^ counter_val_o[31:0];
  assign _055_ = counter_d_t0[63:32] | counter_val_o_t0[63:32];
  assign _059_ = counter_d_t0[31:0] | counter_val_o_t0[31:0];
  assign _056_ = _077_ | _055_;
  assign _060_ = _078_ | _059_;
  assign _030_ = { _008_, _008_, _008_, _008_, _008_, _008_, _008_, _008_, _008_, _008_, _008_, _008_, _008_, _008_, _008_, _008_, _008_, _008_, _008_, _008_, _008_, _008_, _008_, _008_, _008_, _008_, _008_, _008_, _008_, _008_, _008_, _008_ } & counter_d_t0[63:32];
  assign _033_ = { _010_, _010_, _010_, _010_, _010_, _010_, _010_, _010_, _010_, _010_, _010_, _010_, _010_, _010_, _010_, _010_, _010_, _010_, _010_, _010_, _010_, _010_, _010_, _010_, _010_, _010_, _010_, _010_, _010_, _010_, _010_, _010_ } & counter_d_t0[31:0];
  assign _031_ = { _013_, _013_, _013_, _013_, _013_, _013_, _013_, _013_, _013_, _013_, _013_, _013_, _013_, _013_, _013_, _013_, _013_, _013_, _013_, _013_, _013_, _013_, _013_, _013_, _013_, _013_, _013_, _013_, _013_, _013_, _013_, _013_ } & counter_val_o_t0[63:32];
  assign _034_ = { _014_, _014_, _014_, _014_, _014_, _014_, _014_, _014_, _014_, _014_, _014_, _014_, _014_, _014_, _014_, _014_, _014_, _014_, _014_, _014_, _014_, _014_, _014_, _014_, _014_, _014_, _014_, _014_, _014_, _014_, _014_, _014_ } & counter_val_o_t0[31:0];
  assign _032_ = _056_ & { _009_, _009_, _009_, _009_, _009_, _009_, _009_, _009_, _009_, _009_, _009_, _009_, _009_, _009_, _009_, _009_, _009_, _009_, _009_, _009_, _009_, _009_, _009_, _009_, _009_, _009_, _009_, _009_, _009_, _009_, _009_, _009_ };
  assign _035_ = _060_ & { _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_ };
  assign _057_ = _030_ | _031_;
  assign _061_ = _033_ | _034_;
  assign _058_ = _057_ | _032_;
  assign _062_ = _061_ | _035_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) counter_val_o_t0[63:32] <= 32'd0;
    else counter_val_o_t0[63:32] <= _058_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) counter_val_o_t0[31:0] <= 32'd0;
    else counter_val_o_t0[31:0] <= _062_;
  assign _025_ = | { we_t0, counterh_we_i_t0 };
  assign _016_ = ~ { we_t0, counterh_we_i_t0 };
  assign _037_ = { we, counterh_we_i } & _016_;
  assign _038_ = 2'h2 & _016_;
  assign _039_ = 2'h3 & _016_;
  assign _080_ = _037_ == _038_;
  assign _081_ = _037_ == _039_;
  assign _005_ = _080_ & _025_;
  assign _007_ = _081_ & _025_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) counter_val_o[63:32] <= 32'd0;
    else if (_008_) counter_val_o[63:32] <= counter_d[63:32];
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) counter_val_o[31:0] <= 32'd0;
    else if (_010_) counter_val_o[31:0] <= counter_d[31:0];
  assign _024_ = | { we_t0, counter_inc_i_t0 };
  assign _015_ = ~ { we_t0, counter_inc_i_t0 };
  assign _036_ = { we, counter_inc_i } & _015_;
  assign _028_ = ! _036_;
  assign _003_ = _028_ & _024_;
  assign _019_ = ~ { counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i };
  assign _020_ = ~ { we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we };
  assign _021_ = ~ { counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i };
  assign _066_ = { counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0 } | _019_;
  assign _069_ = { we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0 } | _020_;
  assign _072_ = { counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0 } | _021_;
  assign _067_ = { counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0 } | { counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i };
  assign _070_ = { we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0 } | { we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we };
  assign _073_ = { counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0 } | { counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i };
  assign _043_ = 64'h0000000000000000 & _066_;
  assign _046_ = _001_ & _069_;
  assign _049_ = 32'd0 & _072_;
  assign _052_ = counter_val_i_t0 & _072_;
  assign _044_ = counter_upd_t0 & _067_;
  assign _047_ = counter_load_t0 & _070_;
  assign _050_ = counter_val_i_t0 & _073_;
  assign _053_ = 32'd0 & _073_;
  assign _068_ = _043_ | _044_;
  assign _071_ = _046_ | _047_;
  assign _074_ = _049_ | _050_;
  assign _075_ = _052_ | _053_;
  assign _079_ = _000_ ^ counter_load;
  assign _045_ = { counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0 } & counter_upd;
  assign _048_ = { we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0 } & _079_;
  assign _051_ = { counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0 } & counter_val_i;
  assign _001_ = _045_ | _068_;
  assign counter_d_t0 = _048_ | _071_;
  assign counter_load_t0[63:32] = _051_ | _074_;
  assign counter_load_t0[31:0] = _051_ | _075_;
  assign _002_ = | { we, counter_inc_i };
  assign _004_ = { we, counterh_we_i } != 2'h2;
  assign _006_ = { we, counterh_we_i } != 2'h3;
  assign _008_ = & { _004_, _002_ };
  assign _010_ = & { _006_, _002_ };
  assign _017_ = ~ counter_we_i;
  assign _018_ = ~ counterh_we_i;
  assign _040_ = counter_we_i_t0 & _018_;
  assign _041_ = counterh_we_i_t0 & _017_;
  assign _042_ = counter_we_i_t0 & counterh_we_i_t0;
  assign _065_ = _040_ | _041_;
  assign we_t0 = _065_ | _042_;
  assign _026_ = | { _005_, _003_ };
  assign _027_ = | { _007_, _003_ };
  assign _063_ = { _004_, _002_ } | { _005_, _003_ };
  assign _064_ = { _006_, _002_ } | { _007_, _003_ };
  assign _022_ = & _063_;
  assign _023_ = & _064_;
  assign _009_ = _026_ & _022_;
  assign _011_ = _027_ & _023_;
  assign we = counter_we_i | counterh_we_i;
  assign _000_ = counter_inc_i ? counter_upd : 64'hxxxxxxxxxxxxxxxx;
  assign counter_d = we ? counter_load : _000_;
  assign counter_load[63:32] = counterh_we_i ? counter_val_i : 32'hxxxxxxxx;
  assign counter_load[31:0] = counterh_we_i ? 32'hxxxxxxxx : counter_val_i;
endmodule

module paramodauxy_ibex_fetch_fifoNUM_REQS3200000000000000000000000000000010 (clk_i, rst_ni, clear_i, busy_o, in_valid_i, in_addr_i, in_rdata_i, in_err_i, out_valid_o, out_ready_i, out_addr_o, out_addr_next_o, out_rdata_o, out_err_o, out_err_plus2_o, out_valid_o_t0, out_ready_i_t0, out_rdata_o_t0, out_err_plus2_o_t0, out_err_o_t0, out_addr_o_t0
, out_addr_next_o_t0, in_valid_i_t0, in_rdata_i_t0, in_err_i_t0, in_addr_i_t0, clear_i_t0, busy_o_t0);
  wire _000_;
  wire _001_;
  wire _002_;
  wire _003_;
  wire _004_;
  wire _005_;
  wire _006_;
  wire _007_;
  wire _008_;
  wire _009_;
  wire _010_;
  wire _011_;
  wire _012_;
  wire _013_;
  wire _014_;
  wire _015_;
  wire _016_;
  wire _017_;
  wire _018_;
  wire _019_;
  wire _020_;
  wire _021_;
  wire _022_;
  wire _023_;
  wire _024_;
  wire _025_;
  wire _026_;
  wire _027_;
  wire _028_;
  wire _029_;
  wire [30:0] _030_;
  wire [30:0] _031_;
  wire _032_;
  wire _033_;
  wire _034_;
  wire _035_;
  wire [1:0] _036_;
  wire [1:0] _037_;
  wire _038_;
  wire _039_;
  wire _040_;
  wire _041_;
  wire _042_;
  wire _043_;
  wire _044_;
  wire _045_;
  wire _046_;
  wire _047_;
  wire _048_;
  wire _049_;
  wire _050_;
  wire _051_;
  wire _052_;
  wire _053_;
  wire _054_;
  wire [31:0] _055_;
  wire [31:0] _056_;
  wire [31:0] _057_;
  wire [30:0] _058_;
  wire _059_;
  wire [31:0] _060_;
  wire _061_;
  wire _062_;
  wire _063_;
  wire [30:0] _064_;
  wire [30:0] _065_;
  wire _066_;
  wire _067_;
  wire _068_;
  wire _069_;
  wire _070_;
  wire _071_;
  wire _072_;
  wire _073_;
  wire _074_;
  wire _075_;
  wire _076_;
  wire _077_;
  wire _078_;
  wire _079_;
  wire _080_;
  wire _081_;
  wire _082_;
  wire _083_;
  wire _084_;
  wire _085_;
  wire _086_;
  wire _087_;
  wire _088_;
  wire _089_;
  wire _090_;
  wire _091_;
  wire _092_;
  wire _093_;
  wire _094_;
  wire _095_;
  wire _096_;
  wire _097_;
  wire _098_;
  wire _099_;
  wire _100_;
  wire _101_;
  wire _102_;
  wire _103_;
  wire _104_;
  wire _105_;
  wire _106_;
  wire _107_;
  wire _108_;
  wire _109_;
  wire _110_;
  wire _111_;
  wire _112_;
  wire _113_;
  wire _114_;
  wire _115_;
  wire _116_;
  wire _117_;
  wire _118_;
  wire _119_;
  wire _120_;
  wire _121_;
  wire _122_;
  wire _123_;
  wire _124_;
  wire _125_;
  wire _126_;
  wire _127_;
  wire _128_;
  wire _129_;
  wire _130_;
  wire _131_;
  wire _132_;
  wire _133_;
  wire _134_;
  wire _135_;
  wire [31:0] _136_;
  wire [31:0] _137_;
  wire [31:0] _138_;
  wire _139_;
  wire _140_;
  wire _141_;
  wire [31:0] _142_;
  wire [31:0] _143_;
  wire [31:0] _144_;
  wire _145_;
  wire _146_;
  wire _147_;
  wire [31:0] _148_;
  wire [31:0] _149_;
  wire [31:0] _150_;
  wire [30:0] _151_;
  wire [30:0] _152_;
  wire [30:0] _153_;
  wire [1:0] _154_;
  wire [1:0] _155_;
  wire [1:0] _156_;
  wire [1:0] _157_;
  wire _158_;
  wire _159_;
  wire _160_;
  wire _161_;
  wire _162_;
  wire _163_;
  wire _164_;
  wire _165_;
  wire _166_;
  wire _167_;
  wire _168_;
  wire _169_;
  wire _170_;
  wire _171_;
  wire _172_;
  wire _173_;
  wire _174_;
  wire _175_;
  wire _176_;
  wire _177_;
  wire _178_;
  wire _179_;
  wire _180_;
  wire _181_;
  wire _182_;
  wire _183_;
  wire _184_;
  wire _185_;
  wire _186_;
  wire _187_;
  wire _188_;
  wire _189_;
  wire _190_;
  wire _191_;
  wire _192_;
  wire _193_;
  wire _194_;
  wire _195_;
  wire _196_;
  wire _197_;
  wire _198_;
  wire _199_;
  wire [31:0] _200_;
  wire [31:0] _201_;
  wire [31:0] _202_;
  wire [31:0] _203_;
  wire [31:0] _204_;
  wire [31:0] _205_;
  wire _206_;
  wire _207_;
  wire _208_;
  wire [31:0] _209_;
  wire [31:0] _210_;
  wire [31:0] _211_;
  wire _212_;
  wire _213_;
  wire _214_;
  wire _215_;
  wire _216_;
  wire _217_;
  wire _218_;
  wire _219_;
  wire _220_;
  wire _221_;
  wire _222_;
  wire [30:0] _223_;
  wire [30:0] _224_;
  wire [30:0] _225_;
  wire _226_;
  wire _227_;
  wire _228_;
  wire _229_;
  wire _230_;
  wire _231_;
  wire [31:0] _232_;
  wire [31:0] _233_;
  wire [31:0] _234_;
  wire [31:0] _235_;
  wire [31:0] _236_;
  wire [31:0] _237_;
  wire _238_;
  wire _239_;
  wire _240_;
  wire _241_;
  wire _242_;
  wire _243_;
  wire _244_;
  wire [30:0] _245_;
  wire [30:0] _246_;
  wire [30:0] _247_;
  wire _248_;
  wire _249_;
  wire _250_;
  wire _251_;
  wire _252_;
  wire _253_;
  wire _254_;
  wire _255_;
  wire _256_;
  wire _257_;
  wire _258_;
  wire _259_;
  wire _260_;
  wire _261_;
  wire _262_;
  wire _263_;
  wire _264_;
  wire _265_;
  wire _266_;
  wire _267_;
  wire _268_;
  wire _269_;
  wire _270_;
  wire _271_;
  wire _272_;
  wire _273_;
  wire _274_;
  wire [31:0] _275_;
  wire [31:0] _276_;
  wire [31:0] _277_;
  wire [31:0] _278_;
  wire _279_;
  wire _280_;
  wire _281_;
  wire _282_;
  wire [31:0] _283_;
  wire [31:0] _284_;
  wire [31:0] _285_;
  wire [31:0] _286_;
  wire _287_;
  wire _288_;
  wire _289_;
  wire _290_;
  wire [31:0] _291_;
  wire [31:0] _292_;
  wire [31:0] _293_;
  wire [31:0] _294_;
  wire [30:0] _295_;
  wire [30:0] _296_;
  wire [30:0] _297_;
  wire [30:0] _298_;
  wire _299_;
  wire _300_;
  wire _301_;
  wire _302_;
  wire _303_;
  wire _304_;
  wire _305_;
  wire _306_;
  wire _307_;
  wire _308_;
  wire _309_;
  wire _310_;
  wire _311_;
  wire _312_;
  wire _313_;
  wire _314_;
  wire _315_;
  wire _316_;
  wire [31:0] _317_;
  wire [31:0] _318_;
  wire [31:0] _319_;
  wire [31:0] _320_;
  wire [31:0] _321_;
  wire [31:0] _322_;
  wire _323_;
  wire _324_;
  wire _325_;
  wire [31:0] _326_;
  wire [31:0] _327_;
  wire [31:0] _328_;
  wire _329_;
  wire _330_;
  wire _331_;
  wire _332_;
  wire _333_;
  wire [30:0] _334_;
  wire [30:0] _335_;
  wire [30:0] _336_;
  wire _337_;
  wire _338_;
  wire _339_;
  wire _340_;
  wire [31:0] _341_;
  wire [31:0] _342_;
  wire [31:0] _343_;
  wire [31:0] _344_;
  wire _345_;
  wire _346_;
  wire _347_;
  wire _348_;
  wire [30:0] _349_;
  wire _350_;
  wire [31:0] _351_;
  wire _352_;
  wire [31:0] _353_;
  wire _354_;
  wire [31:0] _355_;
  wire [30:0] _356_;
  wire _357_;
  wire _358_;
  wire _359_;
  wire [31:0] _360_;
  wire [31:0] _361_;
  wire _362_;
  wire [31:0] _363_;
  wire _364_;
  wire _365_;
  wire _366_;
  wire [30:0] _367_;
  wire _368_;
  wire _369_;
  wire [31:0] _370_;
  wire _371_;
  wire _372_;
  wire _373_;
  wire [30:0] _374_;
  wire [30:0] _375_;
  wire _376_;
  wire _377_;
  wire _378_;
  wire _379_;
  wire _380_;
  wire _381_;
  wire _382_;
  wire _383_;
  wire _384_;
  wire _385_;
  wire _386_;
  wire _387_;
  wire _388_;
  wire _389_;
  wire _390_;
  wire addr_incr_two;
  wire addr_incr_two_t0;
  wire aligned_is_compressed;
  wire aligned_is_compressed_t0;
  output [1:0] busy_o;
  wire [1:0] busy_o;
  output [1:0] busy_o_t0;
  wire [1:0] busy_o_t0;
  input clear_i;
  wire clear_i;
  input clear_i_t0;
  wire clear_i_t0;
  input clk_i;
  wire clk_i;
  wire [2:0] entry_en;
  wire [2:0] entry_en_t0;
  wire err;
  wire [2:0] err_d;
  wire [2:0] err_d_t0;
  wire err_plus2;
  wire err_plus2_t0;
  reg [2:0] err_q;
  reg [2:0] err_q_t0;
  wire err_t0;
  wire err_unaligned;
  wire err_unaligned_t0;
  input [31:0] in_addr_i;
  wire [31:0] in_addr_i;
  input [31:0] in_addr_i_t0;
  wire [31:0] in_addr_i_t0;
  input in_err_i;
  wire in_err_i;
  input in_err_i_t0;
  wire in_err_i_t0;
  input [31:0] in_rdata_i;
  wire [31:0] in_rdata_i;
  input [31:0] in_rdata_i_t0;
  wire [31:0] in_rdata_i_t0;
  input in_valid_i;
  wire in_valid_i;
  input in_valid_i_t0;
  wire in_valid_i_t0;
  wire [31:1] instr_addr_d;
  wire [31:1] instr_addr_d_t0;
  wire instr_addr_en;
  wire instr_addr_en_t0;
  wire [31:1] instr_addr_next;
  wire [31:1] instr_addr_next_t0;
  reg [31:1] instr_addr_q;
  reg [31:1] instr_addr_q_t0;
  wire [2:0] lowest_free_entry;
  wire [2:0] lowest_free_entry_t0;
  output [31:0] out_addr_next_o;
  wire [31:0] out_addr_next_o;
  output [31:0] out_addr_next_o_t0;
  wire [31:0] out_addr_next_o_t0;
  output [31:0] out_addr_o;
  wire [31:0] out_addr_o;
  output [31:0] out_addr_o_t0;
  wire [31:0] out_addr_o_t0;
  output out_err_o;
  wire out_err_o;
  output out_err_o_t0;
  wire out_err_o_t0;
  output out_err_plus2_o;
  wire out_err_plus2_o;
  output out_err_plus2_o_t0;
  wire out_err_plus2_o_t0;
  output [31:0] out_rdata_o;
  wire [31:0] out_rdata_o;
  output [31:0] out_rdata_o_t0;
  wire [31:0] out_rdata_o_t0;
  input out_ready_i;
  wire out_ready_i;
  input out_ready_i_t0;
  wire out_ready_i_t0;
  output out_valid_o;
  wire out_valid_o;
  output out_valid_o_t0;
  wire out_valid_o_t0;
  wire pop_fifo;
  wire pop_fifo_t0;
  wire [31:0] rdata;
  wire [95:0] rdata_d;
  wire [95:0] rdata_d_t0;
  reg [95:0] rdata_q;
  reg [95:0] rdata_q_t0;
  wire [31:0] rdata_t0;
  wire [31:0] rdata_unaligned;
  wire [31:0] rdata_unaligned_t0;
  input rst_ni;
  wire rst_ni;
  wire unaligned_is_compressed;
  wire unaligned_is_compressed_t0;
  wire valid;
  wire [2:0] valid_d;
  wire [2:0] valid_d_t0;
  wire [2:0] valid_popped;
  wire [2:0] valid_popped_t0;
  wire [2:0] valid_pushed;
  wire [2:0] valid_pushed_t0;
  reg [2:0] valid_q;
  reg [2:0] valid_q_t0;
  wire valid_t0;
  wire valid_unaligned;
  wire valid_unaligned_t0;
  assign instr_addr_next = instr_addr_q + { 29'h00000000, _381_, addr_incr_two };
  assign _002_ = err_q[1] & _054_;
  assign _004_ = valid_q[0] & err_q[0];
  assign _006_ = in_err_i & _385_;
  assign _008_ = err_q[1] & _040_;
  assign _010_ = in_err_i & valid_q[0];
  assign _012_ = _010_ & _040_;
  assign _014_ = valid_q[0] & in_valid_i;
  assign unaligned_is_compressed = _376_ & _380_;
  assign aligned_is_compressed = _378_ & _380_;
  assign _016_ = out_ready_i & out_valid_o;
  assign pop_fifo = _016_ & _389_;
  assign lowest_free_entry[1] = _048_ & valid_q[0];
  assign valid_d[0] = valid_popped[0] & _043_;
  assign valid_d[1] = valid_popped[1] & _043_;
  assign _022_ = valid_pushed[1] & pop_fifo;
  assign _018_ = in_valid_i & lowest_free_entry[0];
  assign _024_ = _018_ & _059_;
  assign _026_ = valid_pushed[2] & pop_fifo;
  assign _020_ = in_valid_i & lowest_free_entry[1];
  assign _028_ = _020_ & _059_;
  assign lowest_free_entry[2] = _053_ & valid_q[1];
  assign valid_d[2] = valid_popped[2] & _043_;
  assign entry_en[2] = in_valid_i & lowest_free_entry[2];
  assign _030_ = ~ instr_addr_q_t0;
  assign _031_ = ~ { 29'h00000000, addr_incr_two_t0, addr_incr_two_t0 };
  assign _064_ = instr_addr_q & _030_;
  assign _065_ = { 29'h00000000, _381_, addr_incr_two } & _031_;
  assign _374_ = _064_ + _065_;
  assign _245_ = instr_addr_q | instr_addr_q_t0;
  assign _246_ = { 29'h00000000, _381_, addr_incr_two } | { 29'h00000000, addr_incr_two_t0, addr_incr_two_t0 };
  assign _375_ = _245_ + _246_;
  assign _349_ = _374_ ^ _375_;
  assign _247_ = _349_ | instr_addr_q_t0;
  assign instr_addr_next_t0 = _247_ | { 29'h00000000, addr_incr_two_t0, addr_incr_two_t0 };
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) valid_q_t0 <= 3'h0;
    else valid_q_t0 <= valid_d_t0;
  assign _066_ = err_q_t0[1] & _054_;
  assign _069_ = valid_q_t0[0] & err_q[0];
  assign _072_ = in_err_i_t0 & _385_;
  assign _075_ = err_q_t0[1] & _040_;
  assign _078_ = in_err_i_t0 & valid_q[0];
  assign _081_ = _011_ & _040_;
  assign _087_ = _377_ & _380_;
  assign _090_ = _379_ & _380_;
  assign _093_ = out_ready_i_t0 & out_valid_o;
  assign _096_ = _017_ & _389_;
  assign _099_ = valid_q_t0[1] & valid_q[0];
  assign _102_ = valid_popped_t0[0] & _043_;
  assign _105_ = valid_popped_t0[1] & _043_;
  assign _108_ = valid_pushed_t0[1] & pop_fifo;
  assign _112_ = _019_ & _059_;
  assign _115_ = valid_pushed_t0[2] & pop_fifo;
  assign _118_ = in_valid_i_t0 & lowest_free_entry[1];
  assign _121_ = _021_ & _059_;
  assign _124_ = valid_q_t0[2] & valid_q[1];
  assign _127_ = valid_popped_t0[2] & _043_;
  assign _130_ = in_valid_i_t0 & lowest_free_entry[2];
  assign _067_ = unaligned_is_compressed_t0 & err_q[1];
  assign _070_ = err_q_t0[0] & valid_q[0];
  assign _073_ = _386_ & in_err_i;
  assign _076_ = err_q_t0[0] & err_q[1];
  assign _079_ = valid_q_t0[0] & in_err_i;
  assign _082_ = err_q_t0[0] & _010_;
  assign _085_ = in_valid_i_t0 & valid_q[0];
  assign _088_ = err_t0 & _376_;
  assign _091_ = err_t0 & _378_;
  assign _094_ = out_valid_o_t0 & out_ready_i;
  assign _097_ = _390_ & _016_;
  assign _100_ = valid_q_t0[0] & _048_;
  assign _103_ = clear_i_t0 & valid_popped[0];
  assign _106_ = clear_i_t0 & valid_popped[1];
  assign _109_ = pop_fifo_t0 & valid_pushed[1];
  assign _084_ = valid_q_t0[0] & in_valid_i;
  assign _113_ = pop_fifo_t0 & _018_;
  assign _119_ = lowest_free_entry_t0[1] & in_valid_i;
  assign _122_ = pop_fifo_t0 & _020_;
  assign _125_ = valid_q_t0[1] & _053_;
  assign _128_ = clear_i_t0 & valid_popped[2];
  assign _131_ = lowest_free_entry_t0[2] & in_valid_i;
  assign _068_ = err_q_t0[1] & unaligned_is_compressed_t0;
  assign _071_ = valid_q_t0[0] & err_q_t0[0];
  assign _074_ = in_err_i_t0 & _386_;
  assign _077_ = err_q_t0[1] & err_q_t0[0];
  assign _080_ = in_err_i_t0 & valid_q_t0[0];
  assign _083_ = _011_ & err_q_t0[0];
  assign _089_ = _377_ & err_t0;
  assign _092_ = _379_ & err_t0;
  assign _095_ = out_ready_i_t0 & out_valid_o_t0;
  assign _098_ = _017_ & _390_;
  assign _101_ = valid_q_t0[1] & valid_q_t0[0];
  assign _104_ = valid_popped_t0[0] & clear_i_t0;
  assign _107_ = valid_popped_t0[1] & clear_i_t0;
  assign _110_ = valid_pushed_t0[1] & pop_fifo_t0;
  assign _114_ = _019_ & pop_fifo_t0;
  assign _117_ = valid_pushed_t0[2] & pop_fifo_t0;
  assign _120_ = in_valid_i_t0 & lowest_free_entry_t0[1];
  assign _123_ = _021_ & pop_fifo_t0;
  assign _126_ = valid_q_t0[2] & valid_q_t0[1];
  assign _129_ = valid_popped_t0[2] & clear_i_t0;
  assign _132_ = in_valid_i_t0 & lowest_free_entry_t0[2];
  assign _248_ = _066_ | _067_;
  assign _249_ = _069_ | _070_;
  assign _250_ = _072_ | _073_;
  assign _251_ = _075_ | _076_;
  assign _252_ = _078_ | _079_;
  assign _253_ = _081_ | _082_;
  assign _254_ = _084_ | _085_;
  assign _255_ = _087_ | _088_;
  assign _256_ = _090_ | _091_;
  assign _257_ = _093_ | _094_;
  assign _258_ = _096_ | _097_;
  assign _259_ = _099_ | _100_;
  assign _260_ = _102_ | _103_;
  assign _261_ = _105_ | _106_;
  assign _262_ = _108_ | _109_;
  assign _263_ = _111_ | _084_;
  assign _264_ = _112_ | _113_;
  assign _265_ = _115_ | _116_;
  assign _266_ = _118_ | _119_;
  assign _267_ = _121_ | _122_;
  assign _268_ = _124_ | _125_;
  assign _269_ = _127_ | _128_;
  assign _270_ = _130_ | _131_;
  assign _003_ = _248_ | _068_;
  assign _005_ = _249_ | _071_;
  assign _007_ = _250_ | _074_;
  assign _009_ = _251_ | _077_;
  assign _011_ = _252_ | _080_;
  assign _013_ = _253_ | _083_;
  assign _015_ = _254_ | _086_;
  assign unaligned_is_compressed_t0 = _255_ | _089_;
  assign aligned_is_compressed_t0 = _256_ | _092_;
  assign _017_ = _257_ | _095_;
  assign pop_fifo_t0 = _258_ | _098_;
  assign lowest_free_entry_t0[1] = _259_ | _101_;
  assign valid_d_t0[0] = _260_ | _104_;
  assign valid_d_t0[1] = _261_ | _107_;
  assign _023_ = _262_ | _110_;
  assign _019_ = _263_ | _086_;
  assign _025_ = _264_ | _114_;
  assign _027_ = _265_ | _117_;
  assign _021_ = _266_ | _120_;
  assign _029_ = _267_ | _123_;
  assign lowest_free_entry_t0[2] = _268_ | _126_;
  assign valid_d_t0[2] = _269_ | _129_;
  assign entry_en_t0[2] = _270_ | _132_;
  assign _352_ = err_d[1] ^ err_q[1];
  assign _353_ = rdata_d[63:32] ^ rdata_q[63:32];
  assign _354_ = err_d[0] ^ err_q[0];
  assign _355_ = rdata_d[31:0] ^ rdata_q[31:0];
  assign _356_ = instr_addr_d ^ instr_addr_q;
  assign _033_ = ~ entry_en[1];
  assign _034_ = ~ entry_en[0];
  assign _035_ = ~ instr_addr_en;
  assign _271_ = in_err_i_t0 | err_q_t0[2];
  assign _275_ = in_rdata_i_t0 | rdata_q_t0[95:64];
  assign _279_ = err_d_t0[1] | err_q_t0[1];
  assign _283_ = rdata_d_t0[63:32] | rdata_q_t0[63:32];
  assign _287_ = err_d_t0[0] | err_q_t0[0];
  assign _291_ = rdata_d_t0[31:0] | rdata_q_t0[31:0];
  assign _295_ = instr_addr_d_t0 | instr_addr_q_t0;
  assign _272_ = _350_ | _271_;
  assign _276_ = _351_ | _275_;
  assign _280_ = _352_ | _279_;
  assign _284_ = _353_ | _283_;
  assign _288_ = _354_ | _287_;
  assign _292_ = _355_ | _291_;
  assign _296_ = _356_ | _295_;
  assign _133_ = entry_en[2] & in_err_i_t0;
  assign _136_ = { entry_en[2], entry_en[2], entry_en[2], entry_en[2], entry_en[2], entry_en[2], entry_en[2], entry_en[2], entry_en[2], entry_en[2], entry_en[2], entry_en[2], entry_en[2], entry_en[2], entry_en[2], entry_en[2], entry_en[2], entry_en[2], entry_en[2], entry_en[2], entry_en[2], entry_en[2], entry_en[2], entry_en[2], entry_en[2], entry_en[2], entry_en[2], entry_en[2], entry_en[2], entry_en[2], entry_en[2], entry_en[2] } & in_rdata_i_t0;
  assign _139_ = entry_en[1] & err_d_t0[1];
  assign _142_ = { entry_en[1], entry_en[1], entry_en[1], entry_en[1], entry_en[1], entry_en[1], entry_en[1], entry_en[1], entry_en[1], entry_en[1], entry_en[1], entry_en[1], entry_en[1], entry_en[1], entry_en[1], entry_en[1], entry_en[1], entry_en[1], entry_en[1], entry_en[1], entry_en[1], entry_en[1], entry_en[1], entry_en[1], entry_en[1], entry_en[1], entry_en[1], entry_en[1], entry_en[1], entry_en[1], entry_en[1], entry_en[1] } & rdata_d_t0[63:32];
  assign _145_ = entry_en[0] & err_d_t0[0];
  assign _148_ = { entry_en[0], entry_en[0], entry_en[0], entry_en[0], entry_en[0], entry_en[0], entry_en[0], entry_en[0], entry_en[0], entry_en[0], entry_en[0], entry_en[0], entry_en[0], entry_en[0], entry_en[0], entry_en[0], entry_en[0], entry_en[0], entry_en[0], entry_en[0], entry_en[0], entry_en[0], entry_en[0], entry_en[0], entry_en[0], entry_en[0], entry_en[0], entry_en[0], entry_en[0], entry_en[0], entry_en[0], entry_en[0] } & rdata_d_t0[31:0];
  assign _151_ = { instr_addr_en, instr_addr_en, instr_addr_en, instr_addr_en, instr_addr_en, instr_addr_en, instr_addr_en, instr_addr_en, instr_addr_en, instr_addr_en, instr_addr_en, instr_addr_en, instr_addr_en, instr_addr_en, instr_addr_en, instr_addr_en, instr_addr_en, instr_addr_en, instr_addr_en, instr_addr_en, instr_addr_en, instr_addr_en, instr_addr_en, instr_addr_en, instr_addr_en, instr_addr_en, instr_addr_en, instr_addr_en, instr_addr_en, instr_addr_en, instr_addr_en } & instr_addr_d_t0;
  assign _134_ = _032_ & err_q_t0[2];
  assign _137_ = { _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_ } & rdata_q_t0[95:64];
  assign _140_ = _033_ & err_q_t0[1];
  assign _143_ = { _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_ } & rdata_q_t0[63:32];
  assign _146_ = _034_ & err_q_t0[0];
  assign _149_ = { _034_, _034_, _034_, _034_, _034_, _034_, _034_, _034_, _034_, _034_, _034_, _034_, _034_, _034_, _034_, _034_, _034_, _034_, _034_, _034_, _034_, _034_, _034_, _034_, _034_, _034_, _034_, _034_, _034_, _034_, _034_, _034_ } & rdata_q_t0[31:0];
  assign _152_ = { _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_ } & instr_addr_q_t0;
  assign _135_ = _272_ & entry_en_t0[2];
  assign _138_ = _276_ & entry_en_t0[2];
  assign _141_ = _280_ & entry_en_t0[1];
  assign _144_ = _284_ & entry_en_t0[1];
  assign _147_ = _288_ & entry_en_t0[0];
  assign _150_ = _292_ & entry_en_t0[0];
  assign _153_ = _296_ & instr_addr_en_t0;
  assign _273_ = _133_ | _134_;
  assign _277_ = _136_ | _137_;
  assign _281_ = _139_ | _140_;
  assign _285_ = _142_ | _143_;
  assign _289_ = _145_ | _146_;
  assign _293_ = _148_ | _149_;
  assign _297_ = _151_ | _152_;
  assign _274_ = _273_ | _135_;
  assign _278_ = _277_ | _138_;
  assign _282_ = _281_ | _141_;
  assign _286_ = _285_ | _144_;
  assign _290_ = _289_ | _147_;
  assign _294_ = _293_ | _150_;
  assign _298_ = _297_ | _153_;
  always_ff @(posedge clk_i)
    err_q_t0[2] <= _274_;
  always_ff @(posedge clk_i)
    rdata_q_t0[95:64] <= _278_;
  always_ff @(posedge clk_i)
    err_q_t0[1] <= _282_;
  always_ff @(posedge clk_i)
    rdata_q_t0[63:32] <= _286_;
  always_ff @(posedge clk_i)
    err_q_t0[0] <= _290_;
  always_ff @(posedge clk_i)
    rdata_q_t0[31:0] <= _294_;
  always_ff @(posedge clk_i)
    instr_addr_q_t0 <= _298_;
  assign _062_ = | rdata_t0[17:16];
  assign _063_ = | rdata_t0[1:0];
  assign _036_ = ~ rdata_t0[17:16];
  assign _037_ = ~ rdata_t0[1:0];
  assign _154_ = rdata[17:16] & _036_;
  assign _156_ = rdata[1:0] & _037_;
  assign _155_ = 2'h3 & _036_;
  assign _157_ = 2'h3 & _037_;
  assign _372_ = _154_ == _155_;
  assign _373_ = _156_ == _157_;
  assign _377_ = _372_ & _062_;
  assign _379_ = _373_ & _063_;
  always_ff @(posedge clk_i)
    if (entry_en[2]) err_q[2] <= in_err_i;
  always_ff @(posedge clk_i)
    if (entry_en[2]) rdata_q[95:64] <= in_rdata_i;
  always_ff @(posedge clk_i)
    if (entry_en[1]) err_q[1] <= err_d[1];
  always_ff @(posedge clk_i)
    if (entry_en[1]) rdata_q[63:32] <= rdata_d[63:32];
  always_ff @(posedge clk_i)
    if (entry_en[0]) err_q[0] <= err_d[0];
  always_ff @(posedge clk_i)
    if (entry_en[0]) rdata_q[31:0] <= rdata_d[31:0];
  always_ff @(posedge clk_i)
    if (instr_addr_en) instr_addr_q <= instr_addr_d;
  assign _054_ = ~ unaligned_is_compressed;
  assign _055_ = ~ { instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1] };
  assign _056_ = ~ { valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0] };
  assign lowest_free_entry[0] = ~ valid_q[0];
  assign _045_ = ~ instr_addr_q[1];
  assign _058_ = ~ { clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i };
  assign _059_ = ~ pop_fifo;
  assign _057_ = ~ { valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1] };
  assign _060_ = ~ { valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2] };
  assign _048_ = ~ valid_q[1];
  assign _053_ = ~ valid_q[2];
  assign _310_ = unaligned_is_compressed_t0 | _054_;
  assign _317_ = { instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1] } | _055_;
  assign _320_ = { valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0] } | _056_;
  assign _323_ = valid_q_t0[0] | lowest_free_entry[0];
  assign _326_ = { valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1] } | _057_;
  assign _329_ = valid_q_t0[1] | _048_;
  assign _313_ = instr_addr_q_t0[1] | _045_;
  assign _334_ = { clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0 } | _058_;
  assign _337_ = pop_fifo_t0 | _059_;
  assign _342_ = { valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2] } | _060_;
  assign _346_ = valid_q_t0[2] | _053_;
  assign _311_ = unaligned_is_compressed_t0 | unaligned_is_compressed;
  assign _318_ = { instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1] } | { instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1] };
  assign _321_ = { valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0] } | { valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0] };
  assign _324_ = valid_q_t0[0] | valid_q[0];
  assign _314_ = instr_addr_q_t0[1] | instr_addr_q[1];
  assign _335_ = { clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0 } | { clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i };
  assign _338_ = pop_fifo_t0 | pop_fifo;
  assign _327_ = { valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1] } | { valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1] };
  assign _343_ = { valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2] } | { valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2] };
  assign _330_ = valid_q_t0[1] | valid_q[1];
  assign _347_ = valid_q_t0[2] | valid_q[2];
  assign _189_ = valid_unaligned_t0 & _310_;
  assign _192_ = valid_t0 & _313_;
  assign _197_ = err_t0 & _313_;
  assign _200_ = rdata_t0 & _317_;
  assign _203_ = in_rdata_i_t0 & _320_;
  assign _206_ = in_err_i_t0 & _323_;
  assign _209_ = { in_rdata_i_t0[15:0], rdata_t0[31:16] } & _326_;
  assign _212_ = _388_ & _329_;
  assign _215_ = _013_ & _329_;
  assign _218_ = _015_ & _329_;
  assign _220_ = aligned_is_compressed_t0 & _313_;
  assign _223_ = instr_addr_next_t0 & _334_;
  assign _226_ = valid_pushed_t0[0] & _337_;
  assign _229_ = valid_pushed_t0[1] & _337_;
  assign _232_ = in_rdata_i_t0 & _326_;
  assign _235_ = in_rdata_i_t0 & _342_;
  assign _238_ = in_err_i_t0 & _329_;
  assign _241_ = in_err_i_t0 & _346_;
  assign _244_ = valid_pushed_t0[2] & _337_;
  assign _190_ = valid_t0 & _311_;
  assign _193_ = _001_ & _314_;
  assign _195_ = err_plus2_t0 & _314_;
  assign _198_ = err_unaligned_t0 & _314_;
  assign _201_ = rdata_unaligned_t0 & _318_;
  assign _204_ = rdata_q_t0[31:0] & _321_;
  assign _207_ = err_q_t0[0] & _324_;
  assign _210_ = { rdata_q_t0[47:32], rdata_t0[31:16] } & _327_;
  assign _213_ = _384_ & _330_;
  assign _216_ = _009_ & _330_;
  assign _221_ = unaligned_is_compressed_t0 & _314_;
  assign _224_ = in_addr_i_t0[31:1] & _335_;
  assign _227_ = valid_pushed_t0[1] & _338_;
  assign _230_ = valid_pushed_t0[2] & _338_;
  assign _233_ = rdata_q_t0[63:32] & _327_;
  assign _236_ = rdata_q_t0[95:64] & _343_;
  assign _239_ = err_q_t0[1] & _330_;
  assign _242_ = err_q_t0[2] & _347_;
  assign _312_ = _189_ | _190_;
  assign _315_ = _192_ | _193_;
  assign _316_ = _197_ | _198_;
  assign _319_ = _200_ | _201_;
  assign _322_ = _203_ | _204_;
  assign _325_ = _206_ | _207_;
  assign _328_ = _209_ | _210_;
  assign _331_ = _212_ | _213_;
  assign _332_ = _215_ | _216_;
  assign _333_ = _220_ | _221_;
  assign _336_ = _223_ | _224_;
  assign _339_ = _226_ | _227_;
  assign _340_ = _229_ | _230_;
  assign _341_ = _232_ | _233_;
  assign _344_ = _235_ | _236_;
  assign _345_ = _238_ | _239_;
  assign _348_ = _241_ | _242_;
  assign _357_ = valid_unaligned ^ valid;
  assign _358_ = valid ^ _000_;
  assign _359_ = err ^ err_unaligned;
  assign _360_ = rdata ^ rdata_unaligned;
  assign _361_ = in_rdata_i ^ rdata_q[31:0];
  assign _362_ = in_err_i ^ err_q[0];
  assign _363_ = { in_rdata_i[15:0], rdata[31:16] } ^ { rdata_q[47:32], rdata[31:16] };
  assign _364_ = _387_ ^ _383_;
  assign _365_ = _012_ ^ _008_;
  assign _366_ = aligned_is_compressed ^ unaligned_is_compressed;
  assign _367_ = instr_addr_next ^ in_addr_i[31:1];
  assign _368_ = valid_pushed[0] ^ valid_pushed[1];
  assign _369_ = valid_pushed[1] ^ valid_pushed[2];
  assign _370_ = in_rdata_i ^ rdata_q[63:32];
  assign _351_ = in_rdata_i ^ rdata_q[95:64];
  assign _371_ = in_err_i ^ err_q[1];
  assign _350_ = in_err_i ^ err_q[2];
  assign _191_ = unaligned_is_compressed_t0 & _357_;
  assign _194_ = instr_addr_q_t0[1] & _358_;
  assign _196_ = instr_addr_q_t0[1] & err_plus2;
  assign _199_ = instr_addr_q_t0[1] & _359_;
  assign _202_ = { instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1] } & _360_;
  assign _205_ = { valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0] } & _361_;
  assign _208_ = valid_q_t0[0] & _362_;
  assign _211_ = { valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1] } & _363_;
  assign _214_ = valid_q_t0[1] & _364_;
  assign _217_ = valid_q_t0[1] & _365_;
  assign _219_ = valid_q_t0[1] & _061_;
  assign _222_ = instr_addr_q_t0[1] & _366_;
  assign _225_ = { clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0 } & _367_;
  assign _228_ = pop_fifo_t0 & _368_;
  assign _231_ = pop_fifo_t0 & _369_;
  assign _234_ = { valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1] } & _370_;
  assign _237_ = { valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2] } & _351_;
  assign _240_ = valid_q_t0[1] & _371_;
  assign _243_ = valid_q_t0[2] & _350_;
  assign _116_ = pop_fifo_t0 & valid_pushed[2];
  assign _001_ = _191_ | _312_;
  assign out_valid_o_t0 = _194_ | _315_;
  assign out_err_plus2_o_t0 = _196_ | _195_;
  assign out_err_o_t0 = _199_ | _316_;
  assign out_rdata_o_t0 = _202_ | _319_;
  assign rdata_t0 = _205_ | _322_;
  assign err_t0 = _208_ | _325_;
  assign rdata_unaligned_t0 = _211_ | _328_;
  assign err_unaligned_t0 = _214_ | _331_;
  assign err_plus2_t0 = _217_ | _332_;
  assign valid_unaligned_t0 = _219_ | _218_;
  assign addr_incr_two_t0 = _222_ | _333_;
  assign instr_addr_d_t0 = _225_ | _336_;
  assign valid_popped_t0[0] = _228_ | _339_;
  assign valid_popped_t0[1] = _231_ | _340_;
  assign rdata_d_t0[31:0] = _234_ | _341_;
  assign rdata_d_t0[63:32] = _237_ | _344_;
  assign err_d_t0[0] = _240_ | _345_;
  assign err_d_t0[1] = _243_ | _348_;
  assign valid_popped_t0[2] = _116_ | _244_;
  assign _061_ = ~ _014_;
  assign _039_ = ~ _002_;
  assign _041_ = ~ _004_;
  assign _043_ = ~ clear_i;
  assign _046_ = ~ _018_;
  assign _047_ = ~ _020_;
  assign _049_ = ~ _022_;
  assign _051_ = ~ _026_;
  assign _038_ = ~ in_valid_i;
  assign _040_ = ~ err_q[0];
  assign _042_ = ~ _006_;
  assign _044_ = ~ _016_;
  assign _050_ = ~ _024_;
  assign _052_ = ~ _028_;
  assign _032_ = ~ entry_en[2];
  assign _158_ = valid_q_t0[0] & _038_;
  assign _159_ = _003_ & _040_;
  assign _162_ = valid_q_t0[0] & unaligned_is_compressed;
  assign _165_ = _005_ & _042_;
  assign _168_ = clear_i_t0 & _044_;
  assign _171_ = aligned_is_compressed_t0 & _045_;
  assign _174_ = _019_ & lowest_free_entry[0];
  assign _177_ = _021_ & _048_;
  assign _180_ = _023_ & _050_;
  assign _183_ = _027_ & _052_;
  assign _186_ = valid_q_t0[2] & _032_;
  assign _111_ = in_valid_i_t0 & lowest_free_entry[0];
  assign _160_ = err_q_t0[0] & _039_;
  assign _163_ = unaligned_is_compressed_t0 & valid_q[0];
  assign _166_ = _007_ & _041_;
  assign _169_ = _017_ & _043_;
  assign _172_ = instr_addr_q_t0[1] & aligned_is_compressed;
  assign _175_ = valid_q_t0[0] & _046_;
  assign _178_ = valid_q_t0[1] & _047_;
  assign _181_ = _025_ & _049_;
  assign _184_ = _029_ & _051_;
  assign _187_ = entry_en_t0[2] & _053_;
  assign _086_ = valid_q_t0[0] & in_valid_i_t0;
  assign _161_ = _003_ & err_q_t0[0];
  assign _164_ = valid_q_t0[0] & unaligned_is_compressed_t0;
  assign _167_ = _005_ & _007_;
  assign _170_ = clear_i_t0 & _017_;
  assign _173_ = aligned_is_compressed_t0 & instr_addr_q_t0[1];
  assign _176_ = _019_ & valid_q_t0[0];
  assign _179_ = _021_ & valid_q_t0[1];
  assign _182_ = _023_ & _025_;
  assign _185_ = _027_ & _029_;
  assign _188_ = valid_q_t0[2] & entry_en_t0[2];
  assign _299_ = _158_ | _111_;
  assign _300_ = _159_ | _160_;
  assign _301_ = _162_ | _163_;
  assign _302_ = _165_ | _166_;
  assign _303_ = _168_ | _169_;
  assign _304_ = _171_ | _172_;
  assign _305_ = _174_ | _175_;
  assign _306_ = _177_ | _178_;
  assign _307_ = _180_ | _181_;
  assign _308_ = _183_ | _184_;
  assign _309_ = _186_ | _187_;
  assign valid_t0 = _299_ | _086_;
  assign _384_ = _300_ | _161_;
  assign _386_ = _301_ | _164_;
  assign _388_ = _302_ | _167_;
  assign instr_addr_en_t0 = _303_ | _170_;
  assign _390_ = _304_ | _173_;
  assign valid_pushed_t0[0] = _305_ | _176_;
  assign valid_pushed_t0[1] = _306_ | _179_;
  assign entry_en_t0[0] = _307_ | _182_;
  assign entry_en_t0[1] = _308_ | _185_;
  assign valid_pushed_t0[2] = _309_ | _188_;
  assign _376_ = rdata[17:16] != 2'h3;
  assign _378_ = rdata[1:0] != 2'h3;
  assign _380_ = ~ err;
  assign _381_ = ~ addr_incr_two;
  assign _382_ = ~ aligned_is_compressed;
  assign valid = valid_q[0] | in_valid_i;
  assign _383_ = _002_ | err_q[0];
  assign _385_ = lowest_free_entry[0] | _054_;
  assign _387_ = _004_ | _006_;
  assign instr_addr_en = clear_i | _016_;
  assign _389_ = _382_ | instr_addr_q[1];
  assign valid_pushed[0] = _018_ | valid_q[0];
  assign valid_pushed[1] = _020_ | valid_q[1];
  assign entry_en[0] = _022_ | _024_;
  assign entry_en[1] = _026_ | _028_;
  assign valid_pushed[2] = valid_q[2] | entry_en[2];
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) valid_q <= 3'h0;
    else valid_q <= valid_d;
  assign _000_ = unaligned_is_compressed ? valid : valid_unaligned;
  assign out_valid_o = instr_addr_q[1] ? _000_ : valid;
  assign out_err_plus2_o = instr_addr_q[1] ? err_plus2 : 1'h0;
  assign out_err_o = instr_addr_q[1] ? err_unaligned : err;
  assign out_rdata_o = instr_addr_q[1] ? rdata_unaligned : rdata;
  assign rdata = valid_q[0] ? rdata_q[31:0] : in_rdata_i;
  assign err = valid_q[0] ? err_q[0] : in_err_i;
  assign rdata_unaligned = valid_q[1] ? { rdata_q[47:32], rdata[31:16] } : { in_rdata_i[15:0], rdata[31:16] };
  assign err_unaligned = valid_q[1] ? _383_ : _387_;
  assign err_plus2 = valid_q[1] ? _008_ : _012_;
  assign valid_unaligned = valid_q[1] ? 1'h1 : _014_;
  assign addr_incr_two = instr_addr_q[1] ? unaligned_is_compressed : aligned_is_compressed;
  assign instr_addr_d = clear_i ? in_addr_i[31:1] : instr_addr_next;
  assign valid_popped[0] = pop_fifo ? valid_pushed[1] : valid_pushed[0];
  assign valid_popped[1] = pop_fifo ? valid_pushed[2] : valid_pushed[1];
  assign rdata_d[31:0] = valid_q[1] ? rdata_q[63:32] : in_rdata_i;
  assign rdata_d[63:32] = valid_q[2] ? rdata_q[95:64] : in_rdata_i;
  assign err_d[0] = valid_q[1] ? err_q[1] : in_err_i;
  assign err_d[1] = valid_q[2] ? err_q[2] : in_err_i;
  assign valid_popped[2] = pop_fifo ? 1'h0 : valid_pushed[2];
  assign busy_o = valid_q[2:1];
  assign busy_o_t0 = valid_q_t0[2:1];
  assign err_d[2] = in_err_i;
  assign err_d_t0[2] = in_err_i_t0;
  assign lowest_free_entry_t0[0] = valid_q_t0[0];
  assign out_addr_next_o = { instr_addr_next, 1'h0 };
  assign out_addr_next_o_t0 = { instr_addr_next_t0, 1'h0 };
  assign out_addr_o = { instr_addr_q, 1'h0 };
  assign out_addr_o_t0 = { instr_addr_q_t0, 1'h0 };
  assign rdata_d[95:64] = in_rdata_i;
  assign rdata_d_t0[95:64] = in_rdata_i_t0;
endmodule

module paramodauxy_ibex_multdiv_fastRV32Ms3200000000000000000000000000000011 (clk_i, rst_ni, mult_en_i, div_en_i, mult_sel_i, div_sel_i, operator_i, signed_mode_i, op_a_i, op_b_i, alu_adder_ext_i, alu_adder_i, equal_to_zero_i, data_ind_timing_i, alu_operand_a_o, alu_operand_b_o, imd_val_q_i, imd_val_d_o, imd_val_we_o, multdiv_ready_id_i, multdiv_result_o
, valid_o, valid_o_t0, data_ind_timing_i_t0, imd_val_d_o_t0, imd_val_q_i_t0, imd_val_we_o_t0, operator_i_t0, alu_adder_ext_i_t0, alu_adder_i_t0, alu_operand_a_o_t0, alu_operand_b_o_t0, div_en_i_t0, div_sel_i_t0, equal_to_zero_i_t0, mult_en_i_t0, mult_sel_i_t0, multdiv_ready_id_i_t0, multdiv_result_o_t0, op_a_i_t0, op_b_i_t0, signed_mode_i_t0
);
  wire _0000_;
  wire _0001_;
  wire [33:0] _0002_;
  wire [33:0] _0003_;
  wire [2:0] _0004_;
  wire [2:0] _0005_;
  wire _0006_;
  wire _0007_;
  wire _0008_;
  wire _0009_;
  wire [33:0] _0010_;
  wire [33:0] _0011_;
  wire [33:0] _0012_;
  wire [33:0] _0013_;
  wire [33:0] _0014_;
  wire [33:0] _0015_;
  wire [34:0] _0016_;
  wire [34:0] _0017_;
  wire _0018_;
  wire _0019_;
  wire _0020_;
  wire _0021_;
  wire _0022_;
  wire _0023_;
  wire _0024_;
  wire _0025_;
  wire _0026_;
  wire _0027_;
  wire _0028_;
  wire _0029_;
  wire [34:0] _0030_;
  wire [34:0] _0031_;
  wire [34:0] _0032_;
  wire _0033_;
  wire _0034_;
  wire _0035_;
  wire _0036_;
  wire _0037_;
  wire [1:0] _0038_;
  wire [1:0] _0039_;
  wire [2:0] _0040_;
  wire _0041_;
  wire _0042_;
  wire _0043_;
  wire _0044_;
  wire [2:0] _0045_;
  wire _0046_;
  wire [33:0] _0047_;
  wire [32:0] _0048_;
  wire [32:0] _0049_;
  wire [32:0] _0050_;
  wire [2:0] _0051_;
  wire [2:0] _0052_;
  wire [2:0] _0053_;
  wire [2:0] _0054_;
  wire [2:0] _0055_;
  wire [2:0] _0056_;
  wire [33:0] _0057_;
  wire [33:0] _0058_;
  wire [33:0] _0059_;
  wire [33:0] _0060_;
  wire [33:0] _0061_;
  wire [31:0] _0062_;
  wire [4:0] _0063_;
  wire [1:0] _0064_;
  wire [1:0] _0065_;
  wire [32:0] _0066_;
  wire [32:0] _0067_;
  wire _0068_;
  wire _0069_;
  wire _0070_;
  wire [33:0] _0071_;
  wire [33:0] _0072_;
  wire [4:0] _0073_;
  wire [32:0] _0074_;
  wire [2:0] _0075_;
  wire [31:0] _0076_;
  wire _0077_;
  wire [33:0] _0078_;
  wire [31:0] _0079_;
  wire [31:0] _0080_;
  wire [32:0] _0081_;
  wire [2:0] _0082_;
  wire [31:0] _0083_;
  wire [31:0] _0084_;
  wire [2:0] _0085_;
  wire [33:0] _0086_;
  wire [33:0] _0087_;
  wire _0088_;
  wire _0089_;
  wire _0090_;
  wire _0091_;
  wire _0092_;
  wire _0093_;
  wire _0094_;
  wire _0095_;
  wire _0096_;
  wire _0097_;
  wire _0098_;
  wire _0099_;
  wire _0100_;
  wire _0101_;
  wire _0102_;
  wire _0103_;
  wire _0104_;
  wire _0105_;
  wire _0106_;
  wire _0107_;
  wire _0108_;
  wire _0109_;
  wire _0110_;
  wire _0111_;
  wire _0112_;
  wire [34:0] _0113_;
  wire [34:0] _0114_;
  wire [34:0] _0115_;
  wire [34:0] _0116_;
  wire _0117_;
  wire _0118_;
  wire _0119_;
  wire _0120_;
  wire _0121_;
  wire _0122_;
  wire _0123_;
  wire _0124_;
  wire _0125_;
  wire _0126_;
  wire _0127_;
  wire _0128_;
  wire _0129_;
  wire _0130_;
  wire _0131_;
  wire _0132_;
  wire _0133_;
  wire _0134_;
  wire [2:0] _0135_;
  wire [2:0] _0136_;
  wire [2:0] _0137_;
  wire [4:0] _0138_;
  wire [4:0] _0139_;
  wire [4:0] _0140_;
  wire _0141_;
  wire _0142_;
  wire _0143_;
  wire [31:0] _0144_;
  wire [31:0] _0145_;
  wire [31:0] _0146_;
  wire [31:0] _0147_;
  wire [31:0] _0148_;
  wire [31:0] _0149_;
  wire _0150_;
  wire _0151_;
  wire _0152_;
  wire [1:0] _0153_;
  wire [1:0] _0154_;
  wire [2:0] _0155_;
  wire _0156_;
  wire _0157_;
  wire _0158_;
  wire _0159_;
  wire _0160_;
  wire _0161_;
  wire [2:0] _0162_;
  wire _0163_;
  wire _0164_;
  wire _0165_;
  wire _0166_;
  wire _0167_;
  wire [33:0] _0168_;
  wire [33:0] _0169_;
  wire [33:0] _0170_;
  wire _0171_;
  wire _0172_;
  wire [33:0] _0173_;
  wire [33:0] _0174_;
  wire [33:0] _0175_;
  wire [33:0] _0176_;
  wire [33:0] _0177_;
  wire [32:0] _0178_;
  wire [32:0] _0179_;
  wire [32:0] _0180_;
  wire [32:0] _0181_;
  wire [32:0] _0182_;
  wire [32:0] _0183_;
  wire [32:0] _0184_;
  wire [32:0] _0185_;
  wire [32:0] _0186_;
  wire [2:0] _0187_;
  wire [2:0] _0188_;
  wire [2:0] _0189_;
  wire [2:0] _0190_;
  wire [2:0] _0191_;
  wire [2:0] _0192_;
  wire [2:0] _0193_;
  wire [2:0] _0194_;
  wire [2:0] _0195_;
  wire [2:0] _0196_;
  wire [2:0] _0197_;
  wire [2:0] _0198_;
  wire [2:0] _0199_;
  wire [2:0] _0200_;
  wire [2:0] _0201_;
  wire [2:0] _0202_;
  wire [2:0] _0203_;
  wire [2:0] _0204_;
  wire [33:0] _0205_;
  wire [33:0] _0206_;
  wire [33:0] _0207_;
  wire [33:0] _0208_;
  wire [33:0] _0209_;
  wire [33:0] _0210_;
  wire [33:0] _0211_;
  wire [33:0] _0212_;
  wire [33:0] _0213_;
  wire [33:0] _0214_;
  wire [33:0] _0215_;
  wire [33:0] _0216_;
  wire [33:0] _0217_;
  wire [33:0] _0218_;
  wire [33:0] _0219_;
  wire [31:0] _0220_;
  wire [31:0] _0221_;
  wire [31:0] _0222_;
  wire [4:0] _0223_;
  wire [4:0] _0224_;
  wire [1:0] _0225_;
  wire [1:0] _0226_;
  wire _0227_;
  wire _0228_;
  wire _0229_;
  wire [1:0] _0230_;
  wire _0231_;
  wire _0232_;
  wire _0233_;
  wire [32:0] _0234_;
  wire [32:0] _0235_;
  wire [32:0] _0236_;
  wire _0237_;
  wire _0238_;
  wire _0239_;
  wire _0240_;
  wire _0241_;
  wire [33:0] _0242_;
  wire [33:0] _0243_;
  wire [33:0] _0244_;
  wire _0245_;
  wire _0246_;
  wire [33:0] _0247_;
  wire [33:0] _0248_;
  wire [33:0] _0249_;
  wire [33:0] _0250_;
  wire [33:0] _0251_;
  wire [33:0] _0252_;
  wire [33:0] _0253_;
  wire [33:0] _0254_;
  wire [33:0] _0255_;
  wire [4:0] _0256_;
  wire [4:0] _0257_;
  wire [4:0] _0258_;
  wire [32:0] _0259_;
  wire [32:0] _0260_;
  wire [32:0] _0261_;
  wire [2:0] _0262_;
  wire [2:0] _0263_;
  wire [2:0] _0264_;
  wire _0265_;
  wire _0266_;
  wire [2:0] _0267_;
  wire [2:0] _0268_;
  wire [2:0] _0269_;
  wire [31:0] _0270_;
  wire [31:0] _0271_;
  wire [31:0] _0272_;
  wire [2:0] _0273_;
  wire _0274_;
  wire _0275_;
  wire _0276_;
  wire [33:0] _0277_;
  wire [33:0] _0278_;
  wire [33:0] _0279_;
  wire [31:0] _0280_;
  wire [31:0] _0281_;
  wire [31:0] _0282_;
  wire [31:0] _0283_;
  wire [31:0] _0284_;
  wire [31:0] _0285_;
  wire [32:0] _0286_;
  wire [32:0] _0287_;
  wire [32:0] _0288_;
  wire [2:0] _0289_;
  wire [2:0] _0290_;
  wire [2:0] _0291_;
  wire [31:0] _0292_;
  wire [31:0] _0293_;
  wire [31:0] _0294_;
  wire [31:0] _0295_;
  wire [31:0] _0296_;
  wire [31:0] _0297_;
  wire [2:0] _0298_;
  wire [2:0] _0299_;
  wire [2:0] _0300_;
  wire [33:0] _0301_;
  wire [33:0] _0302_;
  wire [33:0] _0303_;
  wire [33:0] _0304_;
  wire [33:0] _0305_;
  wire [33:0] _0306_;
  wire _0307_;
  wire _0308_;
  wire _0309_;
  wire _0310_;
  wire [34:0] _0311_;
  wire [34:0] _0312_;
  wire [34:0] _0313_;
  wire [34:0] _0314_;
  wire _0315_;
  wire _0316_;
  wire _0317_;
  wire _0318_;
  wire _0319_;
  wire _0320_;
  wire [2:0] _0321_;
  wire [2:0] _0322_;
  wire [2:0] _0323_;
  wire [2:0] _0324_;
  wire [4:0] _0325_;
  wire [4:0] _0326_;
  wire [4:0] _0327_;
  wire [4:0] _0328_;
  wire _0329_;
  wire _0330_;
  wire _0331_;
  wire _0332_;
  wire [31:0] _0333_;
  wire [31:0] _0334_;
  wire [31:0] _0335_;
  wire [31:0] _0336_;
  wire [31:0] _0337_;
  wire [31:0] _0338_;
  wire [31:0] _0339_;
  wire [31:0] _0340_;
  wire _0341_;
  wire _0342_;
  wire _0343_;
  wire _0344_;
  wire [1:0] _0345_;
  wire [1:0] _0346_;
  wire [2:0] _0347_;
  wire _0348_;
  wire _0349_;
  wire _0350_;
  wire _0351_;
  wire _0352_;
  wire [33:0] _0353_;
  wire [33:0] _0354_;
  wire [33:0] _0355_;
  wire [33:0] _0356_;
  wire [33:0] _0357_;
  wire [32:0] _0358_;
  wire [32:0] _0359_;
  wire [32:0] _0360_;
  wire [32:0] _0361_;
  wire [32:0] _0362_;
  wire [32:0] _0363_;
  wire [32:0] _0364_;
  wire [32:0] _0365_;
  wire [32:0] _0366_;
  wire [2:0] _0367_;
  wire [2:0] _0368_;
  wire [2:0] _0369_;
  wire [2:0] _0370_;
  wire [2:0] _0371_;
  wire [2:0] _0372_;
  wire [2:0] _0373_;
  wire [2:0] _0374_;
  wire [2:0] _0375_;
  wire [2:0] _0376_;
  wire [2:0] _0377_;
  wire [2:0] _0378_;
  wire [2:0] _0379_;
  wire [2:0] _0380_;
  wire [2:0] _0381_;
  wire [2:0] _0382_;
  wire [2:0] _0383_;
  wire [2:0] _0384_;
  wire [33:0] _0385_;
  wire [33:0] _0386_;
  wire [33:0] _0387_;
  wire [33:0] _0388_;
  wire [33:0] _0389_;
  wire [33:0] _0390_;
  wire [33:0] _0391_;
  wire [33:0] _0392_;
  wire [33:0] _0393_;
  wire [33:0] _0394_;
  wire [33:0] _0395_;
  wire [33:0] _0396_;
  wire [33:0] _0397_;
  wire [33:0] _0398_;
  wire [33:0] _0399_;
  wire [31:0] _0400_;
  wire [31:0] _0401_;
  wire [31:0] _0402_;
  wire _0403_;
  wire _0404_;
  wire [32:0] _0405_;
  wire _0406_;
  wire _0407_;
  wire [33:0] _0408_;
  wire [33:0] _0409_;
  wire [33:0] _0410_;
  wire [33:0] _0411_;
  wire [33:0] _0412_;
  wire [33:0] _0413_;
  wire [33:0] _0414_;
  wire [33:0] _0415_;
  wire [4:0] _0416_;
  wire [4:0] _0417_;
  wire [4:0] _0418_;
  wire [32:0] _0419_;
  wire [32:0] _0420_;
  wire [32:0] _0421_;
  wire _0422_;
  wire [31:0] _0423_;
  wire [31:0] _0424_;
  wire [31:0] _0425_;
  wire _0426_;
  wire _0427_;
  wire _0428_;
  wire [4:0] _0429_;
  wire [4:0] _0430_;
  wire [33:0] _0431_;
  wire [33:0] _0432_;
  wire [33:0] _0433_;
  wire [31:0] _0434_;
  wire [31:0] _0435_;
  wire [31:0] _0436_;
  wire [31:0] _0437_;
  wire [31:0] _0438_;
  wire [31:0] _0439_;
  wire [32:0] _0440_;
  wire [32:0] _0441_;
  wire [32:0] _0442_;
  wire [2:0] _0443_;
  wire [2:0] _0444_;
  wire [2:0] _0445_;
  wire [31:0] _0446_;
  wire [31:0] _0447_;
  wire [31:0] _0448_;
  wire [31:0] _0449_;
  wire [31:0] _0450_;
  wire [31:0] _0451_;
  wire [2:0] _0452_;
  wire [2:0] _0453_;
  wire [2:0] _0454_;
  wire [33:0] _0455_;
  wire [33:0] _0456_;
  wire [33:0] _0457_;
  wire [33:0] _0458_;
  wire [33:0] _0459_;
  wire [33:0] _0460_;
  wire [34:0] _0461_;
  wire [34:0] _0462_;
  wire [2:0] _0463_;
  wire [4:0] _0464_;
  wire _0465_;
  wire [31:0] _0466_;
  wire [31:0] _0467_;
  wire _0468_;
  wire _0469_;
  wire [33:0] _0470_;
  wire [33:0] _0471_;
  wire [32:0] _0472_;
  wire [32:0] _0473_;
  wire [32:0] _0474_;
  wire [2:0] _0475_;
  wire [2:0] _0476_;
  wire [2:0] _0477_;
  wire [2:0] _0478_;
  wire [33:0] _0479_;
  wire [33:0] _0480_;
  wire [33:0] _0481_;
  wire [33:0] _0482_;
  wire [33:0] _0483_;
  wire [33:0] _0484_;
  wire _0485_;
  wire [33:0] _0486_;
  wire [33:0] _0487_;
  wire [33:0] _0488_;
  wire [4:0] _0489_;
  wire [32:0] _0490_;
  wire [31:0] _0491_;
  wire _0492_;
  wire [4:0] _0493_;
  wire [33:0] _0494_;
  wire [31:0] _0495_;
  wire [31:0] _0496_;
  wire [32:0] _0497_;
  wire [31:0] _0498_;
  wire [31:0] _0499_;
  wire [33:0] _0500_;
  wire _0501_;
  wire _0502_;
  wire _0503_;
  wire _0504_;
  wire _0505_;
  wire _0506_;
  wire _0507_;
  wire _0508_;
  wire [34:0] _0509_;
  wire [34:0] _0510_;
  wire [34:0] _0511_;
  wire [34:0] _0512_;
  wire [4:0] _0513_;
  wire [4:0] _0514_;
  wire [32:0] _0515_;
  wire [32:0] _0516_;
  wire [32:0] _0517_;
  wire [32:0] _0518_;
  wire [2:0] _0519_;
  wire [2:0] _0520_;
  wire [2:0] _0521_;
  wire [2:0] _0522_;
  wire [2:0] _0523_;
  wire [2:0] _0524_;
  wire [2:0] _0525_;
  wire [2:0] _0526_;
  wire [2:0] _0527_;
  wire [2:0] _0528_;
  wire [33:0] _0529_;
  wire [33:0] _0530_;
  wire [33:0] _0531_;
  wire [33:0] _0532_;
  wire [33:0] _0533_;
  wire [33:0] _0534_;
  wire [33:0] _0535_;
  wire [33:0] _0536_;
  wire _0537_;
  wire [31:0] _0538_;
  wire _0539_;
  wire _0540_;
  wire _0541_;
  wire _0542_;
  wire _0543_;
  wire _0544_;
  wire _0545_;
  wire _0546_;
  wire _0547_;
  wire _0548_;
  wire _0549_;
  wire _0550_;
  wire [31:0] _0551_;
  wire [31:0] _0552_;
  wire [31:0] _0553_;
  wire [31:0] _0554_;
  wire [32:0] _0555_;
  wire [32:0] _0556_;
  wire _0557_;
  wire _0558_;
  wire _0559_;
  wire _0560_;
  wire _0561_;
  wire _0562_;
  wire _0563_;
  wire _0564_;
  wire _0565_;
  wire _0566_;
  wire _0567_;
  wire _0568_;
  wire _0569_;
  wire _0570_;
  wire _0571_;
  wire [4:0] _0572_;
  wire [31:0] _0573_;
  wire [31:0] _0574_;
  wire [31:0] _0575_;
  wire [31:0] _0576_;
  wire [2:0] _0577_;
  wire [2:0] _0578_;
  wire [33:0] _0579_;
  wire [33:0] _0580_;
  wire [33:0] _0581_;
  wire [33:0] _0582_;
  wire _0583_;
  wire _0584_;
  wire _0585_;
  wire _0586_;
  wire [33:0] accum;
  wire [33:0] accum_t0;
  input [33:0] alu_adder_ext_i;
  wire [33:0] alu_adder_ext_i;
  input [33:0] alu_adder_ext_i_t0;
  wire [33:0] alu_adder_ext_i_t0;
  input [31:0] alu_adder_i;
  wire [31:0] alu_adder_i;
  input [31:0] alu_adder_i_t0;
  wire [31:0] alu_adder_i_t0;
  output [32:0] alu_operand_a_o;
  wire [32:0] alu_operand_a_o;
  output [32:0] alu_operand_a_o_t0;
  wire [32:0] alu_operand_a_o_t0;
  output [32:0] alu_operand_b_o;
  wire [32:0] alu_operand_b_o;
  output [32:0] alu_operand_b_o_t0;
  wire [32:0] alu_operand_b_o_t0;
  input clk_i;
  wire clk_i;
  input data_ind_timing_i;
  wire data_ind_timing_i;
  input data_ind_timing_i_t0;
  wire data_ind_timing_i_t0;
  reg div_by_zero_q;
  reg div_by_zero_q_t0;
  wire div_change_sign;
  wire div_change_sign_t0;
  wire [4:0] div_counter_d;
  wire [4:0] div_counter_d_t0;
  reg [4:0] div_counter_q;
  reg [4:0] div_counter_q_t0;
  input div_en_i;
  wire div_en_i;
  input div_en_i_t0;
  wire div_en_i_t0;
  wire div_en_internal;
  wire div_en_internal_t0;
  wire div_hold;
  wire div_hold_t0;
  input div_sel_i;
  wire div_sel_i;
  input div_sel_i_t0;
  wire div_sel_i_t0;
  wire div_sign_a;
  wire div_sign_a_t0;
  wire div_sign_b;
  wire div_sign_b_t0;
  wire div_valid;
  wire div_valid_t0;
  input equal_to_zero_i;
  wire equal_to_zero_i;
  input equal_to_zero_i_t0;
  wire equal_to_zero_i_t0;
  wire [33:0] \gen_mult_single_cycle.mult1_res ;
  wire [33:0] \gen_mult_single_cycle.mult2_res ;
  wire [15:0] \gen_mult_single_cycle.mult3_op_b ;
  wire [33:0] \gen_mult_single_cycle.mult3_res ;
  wire \gen_mult_single_cycle.mult3_sign_b ;
  wire \gen_mult_single_cycle.mult_state_d ;
  wire \gen_mult_single_cycle.mult_state_d_t0 ;
  reg \gen_mult_single_cycle.mult_state_q ;
  reg \gen_mult_single_cycle.mult_state_q_t0 ;
  wire [33:0] \gen_mult_single_cycle.summand1 ;
  wire [33:0] \gen_mult_single_cycle.summand1_t0 ;
  wire [33:0] \gen_mult_single_cycle.summand2 ;
  wire [33:0] \gen_mult_single_cycle.summand2_t0 ;
  output [67:0] imd_val_d_o;
  wire [67:0] imd_val_d_o;
  output [67:0] imd_val_d_o_t0;
  wire [67:0] imd_val_d_o_t0;
  input [67:0] imd_val_q_i;
  wire [67:0] imd_val_q_i;
  input [67:0] imd_val_q_i_t0;
  wire [67:0] imd_val_q_i_t0;
  output [1:0] imd_val_we_o;
  wire [1:0] imd_val_we_o;
  output [1:0] imd_val_we_o_t0;
  wire [1:0] imd_val_we_o_t0;
  wire is_greater_equal;
  wire is_greater_equal_t0;
  wire [33:0] mac_res_d;
  wire [33:0] mac_res_d_t0;
  wire [34:0] mac_res_ext;
  wire [34:0] mac_res_ext_t0;
  wire [2:0] md_state_d;
  wire [2:0] md_state_d_t0;
  reg [2:0] md_state_q;
  reg [2:0] md_state_q_t0;
  input mult_en_i;
  wire mult_en_i;
  input mult_en_i_t0;
  wire mult_en_i_t0;
  wire mult_en_internal;
  wire mult_en_internal_t0;
  wire mult_hold;
  wire mult_hold_t0;
  input mult_sel_i;
  wire mult_sel_i;
  input mult_sel_i_t0;
  wire mult_sel_i_t0;
  wire mult_valid;
  wire mult_valid_t0;
  wire multdiv_en;
  wire multdiv_en_t0;
  input multdiv_ready_id_i;
  wire multdiv_ready_id_i;
  input multdiv_ready_id_i_t0;
  wire multdiv_ready_id_i_t0;
  output [31:0] multdiv_result_o;
  wire [31:0] multdiv_result_o;
  output [31:0] multdiv_result_o_t0;
  wire [31:0] multdiv_result_o_t0;
  wire [32:0] next_quotient;
  wire [32:0] next_quotient_t0;
  wire [31:0] next_remainder;
  wire [31:0] next_remainder_t0;
  wire [31:0] one_shift;
  wire [31:0] one_shift_t0;
  input [31:0] op_a_i;
  wire [31:0] op_a_i;
  input [31:0] op_a_i_t0;
  wire [31:0] op_a_i_t0;
  input [31:0] op_b_i;
  wire [31:0] op_b_i;
  input [31:0] op_b_i_t0;
  wire [31:0] op_b_i_t0;
  wire [31:0] op_denominator_d;
  wire [31:0] op_denominator_d_t0;
  reg [31:0] op_numerator_q;
  reg [31:0] op_numerator_q_t0;
  wire [31:0] op_quotient_d;
  wire [31:0] op_quotient_d_t0;
  reg [31:0] op_quotient_q;
  reg [31:0] op_quotient_q_t0;
  wire [33:0] op_remainder_d;
  wire [33:0] op_remainder_d_t0;
  input [1:0] operator_i;
  wire [1:0] operator_i;
  input [1:0] operator_i_t0;
  wire [1:0] operator_i_t0;
  input rst_ni;
  wire rst_ni;
  input [1:0] signed_mode_i;
  wire [1:0] signed_mode_i;
  input [1:0] signed_mode_i_t0;
  wire [1:0] signed_mode_i_t0;
  wire signed_mult;
  wire signed_mult_t0;
  output valid_o;
  wire valid_o;
  output valid_o_t0;
  wire valid_o_t0;
  assign _0016_ = $signed({ \gen_mult_single_cycle.summand1 [33], \gen_mult_single_cycle.summand1  }) + $signed({ \gen_mult_single_cycle.summand2 [33], \gen_mult_single_cycle.summand2  });
  assign mac_res_ext = $signed(_0016_) + $signed({ \gen_mult_single_cycle.mult3_res [33], \gen_mult_single_cycle.mult3_res  });
  assign mult_en_internal = mult_en_i & _0548_;
  assign div_en_internal = div_en_i & _0549_;
  assign div_sign_a = signed_mode_i[0] & op_a_i[31];
  assign div_sign_b = signed_mode_i[1] & op_b_i[31];
  assign accum[33] = signed_mult & imd_val_q_i[67];
  assign div_change_sign = _0585_ & _0550_;
  assign _0030_ = ~ { \gen_mult_single_cycle.summand1_t0 [33], \gen_mult_single_cycle.summand1_t0  };
  assign _0032_ = ~ _0017_;
  assign _0031_ = ~ { \gen_mult_single_cycle.summand2_t0 [33], \gen_mult_single_cycle.summand2_t0  };
  assign _0113_ = { \gen_mult_single_cycle.summand1 [33], \gen_mult_single_cycle.summand1  } & _0030_;
  assign _0115_ = _0016_ & _0032_;
  assign _0114_ = { \gen_mult_single_cycle.summand2 [33], \gen_mult_single_cycle.summand2  } & _0031_;
  assign _0116_ = { \gen_mult_single_cycle.mult3_res [33], \gen_mult_single_cycle.mult3_res  } & 35'h7ffffffff;
  assign _0509_ = _0113_ + _0114_;
  assign _0511_ = _0115_ + _0116_;
  assign _0311_ = { \gen_mult_single_cycle.summand1 [33], \gen_mult_single_cycle.summand1  } | { \gen_mult_single_cycle.summand1_t0 [33], \gen_mult_single_cycle.summand1_t0  };
  assign _0314_ = _0016_ | _0017_;
  assign _0312_ = { \gen_mult_single_cycle.summand2 [33], \gen_mult_single_cycle.summand2  } | { \gen_mult_single_cycle.summand2_t0 [33], \gen_mult_single_cycle.summand2_t0  };
  assign _0510_ = _0311_ + _0312_;
  assign _0512_ = _0314_ + { \gen_mult_single_cycle.mult3_res [33], \gen_mult_single_cycle.mult3_res  };
  assign _0461_ = _0509_ ^ _0510_;
  assign _0462_ = _0511_ ^ _0512_;
  assign _0313_ = _0461_ | { \gen_mult_single_cycle.summand1_t0 [33], \gen_mult_single_cycle.summand1_t0  };
  assign mac_res_ext_t0 = _0462_ | _0017_;
  assign _0017_ = _0313_ | { \gen_mult_single_cycle.summand2_t0 [33], \gen_mult_single_cycle.summand2_t0  };
  assign _0035_ = ~ _0020_;
  assign _0036_ = ~ _0022_;
  assign _0037_ = ~ _0024_;
  assign _0463_ = md_state_d ^ md_state_q;
  assign _0464_ = div_counter_d ^ div_counter_q;
  assign _0465_ = \gen_mult_single_cycle.mult_state_d  ^ \gen_mult_single_cycle.mult_state_q ;
  assign _0466_ = op_quotient_d ^ op_quotient_q;
  assign _0467_ = _0573_ ^ op_numerator_q;
  assign _0468_ = equal_to_zero_i ^ div_by_zero_q;
  assign _0321_ = md_state_d_t0 | md_state_q_t0;
  assign _0325_ = div_counter_d_t0 | div_counter_q_t0;
  assign _0329_ = \gen_mult_single_cycle.mult_state_d_t0  | \gen_mult_single_cycle.mult_state_q_t0 ;
  assign _0333_ = op_quotient_d_t0 | op_quotient_q_t0;
  assign _0337_ = _0574_ | op_numerator_q_t0;
  assign _0341_ = equal_to_zero_i_t0 | div_by_zero_q_t0;
  assign _0322_ = _0463_ | _0321_;
  assign _0326_ = _0464_ | _0325_;
  assign _0330_ = _0465_ | _0329_;
  assign _0334_ = _0466_ | _0333_;
  assign _0338_ = _0467_ | _0337_;
  assign _0342_ = _0468_ | _0341_;
  assign _0135_ = { div_en_internal, div_en_internal, div_en_internal } & md_state_d_t0;
  assign _0138_ = { div_en_internal, div_en_internal, div_en_internal, div_en_internal, div_en_internal } & div_counter_d_t0;
  assign _0141_ = mult_en_internal & \gen_mult_single_cycle.mult_state_d_t0 ;
  assign _0144_ = { _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_ } & op_quotient_d_t0;
  assign _0147_ = { _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_ } & _0574_;
  assign _0150_ = _0024_ & equal_to_zero_i_t0;
  assign _0136_ = { _0033_, _0033_, _0033_ } & md_state_q_t0;
  assign _0139_ = { _0033_, _0033_, _0033_, _0033_, _0033_ } & div_counter_q_t0;
  assign _0142_ = _0034_ & \gen_mult_single_cycle.mult_state_q_t0 ;
  assign _0145_ = { _0035_, _0035_, _0035_, _0035_, _0035_, _0035_, _0035_, _0035_, _0035_, _0035_, _0035_, _0035_, _0035_, _0035_, _0035_, _0035_, _0035_, _0035_, _0035_, _0035_, _0035_, _0035_, _0035_, _0035_, _0035_, _0035_, _0035_, _0035_, _0035_, _0035_, _0035_, _0035_ } & op_quotient_q_t0;
  assign _0148_ = { _0036_, _0036_, _0036_, _0036_, _0036_, _0036_, _0036_, _0036_, _0036_, _0036_, _0036_, _0036_, _0036_, _0036_, _0036_, _0036_, _0036_, _0036_, _0036_, _0036_, _0036_, _0036_, _0036_, _0036_, _0036_, _0036_, _0036_, _0036_, _0036_, _0036_, _0036_, _0036_ } & op_numerator_q_t0;
  assign _0151_ = _0037_ & div_by_zero_q_t0;
  assign _0137_ = _0322_ & { div_en_internal_t0, div_en_internal_t0, div_en_internal_t0 };
  assign _0140_ = _0326_ & { div_en_internal_t0, div_en_internal_t0, div_en_internal_t0, div_en_internal_t0, div_en_internal_t0 };
  assign _0143_ = _0330_ & mult_en_internal_t0;
  assign _0146_ = _0334_ & { _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_ };
  assign _0149_ = _0338_ & { _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_ };
  assign _0152_ = _0342_ & _0025_;
  assign _0323_ = _0135_ | _0136_;
  assign _0327_ = _0138_ | _0139_;
  assign _0331_ = _0141_ | _0142_;
  assign _0335_ = _0144_ | _0145_;
  assign _0339_ = _0147_ | _0148_;
  assign _0343_ = _0150_ | _0151_;
  assign _0324_ = _0323_ | _0137_;
  assign _0328_ = _0327_ | _0140_;
  assign _0332_ = _0331_ | _0143_;
  assign _0336_ = _0335_ | _0146_;
  assign _0340_ = _0339_ | _0149_;
  assign _0344_ = _0343_ | _0152_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) md_state_q_t0 <= 3'h0;
    else md_state_q_t0 <= _0324_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) div_counter_q_t0 <= 5'h00;
    else div_counter_q_t0 <= _0328_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) \gen_mult_single_cycle.mult_state_q_t0  <= 1'h0;
    else \gen_mult_single_cycle.mult_state_q_t0  <= _0332_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) op_quotient_q_t0 <= 32'd0;
    else op_quotient_q_t0 <= _0336_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) op_numerator_q_t0 <= 32'd0;
    else op_numerator_q_t0 <= _0340_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) div_by_zero_q_t0 <= 1'h0;
    else div_by_zero_q_t0 <= _0344_;
  assign _0117_ = mult_en_i_t0 & _0548_;
  assign _0120_ = div_en_i_t0 & _0549_;
  assign _0123_ = signed_mode_i_t0[0] & op_a_i[31];
  assign _0126_ = signed_mode_i_t0[1] & op_b_i[31];
  assign _0129_ = signed_mult_t0 & imd_val_q_i[67];
  assign _0132_ = _0586_ & _0550_;
  assign _0118_ = mult_hold_t0 & mult_en_i;
  assign _0121_ = div_hold_t0 & div_en_i;
  assign _0124_ = op_a_i_t0[31] & signed_mode_i[0];
  assign _0127_ = op_b_i_t0[31] & signed_mode_i[1];
  assign _0130_ = imd_val_q_i_t0[67] & signed_mult;
  assign _0133_ = div_by_zero_q_t0 & _0585_;
  assign _0119_ = mult_en_i_t0 & mult_hold_t0;
  assign _0122_ = div_en_i_t0 & div_hold_t0;
  assign _0125_ = signed_mode_i_t0[0] & op_a_i_t0[31];
  assign _0128_ = signed_mode_i_t0[1] & op_b_i_t0[31];
  assign _0131_ = signed_mult_t0 & imd_val_q_i_t0[67];
  assign _0134_ = _0586_ & div_by_zero_q_t0;
  assign _0315_ = _0117_ | _0118_;
  assign _0316_ = _0120_ | _0121_;
  assign _0317_ = _0123_ | _0124_;
  assign _0318_ = _0126_ | _0127_;
  assign _0319_ = _0129_ | _0130_;
  assign _0320_ = _0132_ | _0133_;
  assign mult_en_internal_t0 = _0315_ | _0119_;
  assign div_en_internal_t0 = _0316_ | _0122_;
  assign div_sign_a_t0 = _0317_ | _0125_;
  assign div_sign_b_t0 = _0318_ | _0128_;
  assign accum_t0[33] = _0319_ | _0131_;
  assign div_change_sign_t0 = _0320_ | _0134_;
  assign _0104_ = | md_state_q_t0;
  assign _0063_ = ~ div_counter_q_t0;
  assign _0064_ = ~ operator_i_t0;
  assign _0075_ = ~ md_state_q_t0;
  assign _0223_ = div_counter_q & _0063_;
  assign _0225_ = operator_i & _0064_;
  assign _0262_ = md_state_q & _0075_;
  assign _0224_ = 5'h01 & _0063_;
  assign _0226_ = 2'h2 & _0064_;
  assign _0263_ = 3'h5 & _0075_;
  assign _0264_ = 3'h4 & _0075_;
  assign _0267_ = 3'h6 & _0075_;
  assign _0268_ = 3'h3 & _0075_;
  assign _0269_ = 3'h1 & _0075_;
  assign _0273_ = 3'h2 & _0075_;
  assign _0501_ = _0223_ == _0224_;
  assign _0502_ = _0225_ == _0226_;
  assign _0503_ = _0262_ == _0263_;
  assign _0504_ = _0262_ == _0264_;
  assign _0505_ = _0262_ == _0267_;
  assign _0506_ = _0262_ == _0268_;
  assign _0507_ = _0262_ == _0269_;
  assign _0508_ = _0262_ == _0273_;
  assign _0543_ = _0501_ & _0101_;
  assign _0541_ = _0502_ & _0102_;
  assign _0558_ = _0503_ & _0104_;
  assign _0560_ = _0504_ & _0104_;
  assign div_valid_t0 = _0505_ & _0104_;
  assign _0568_ = _0506_ & _0104_;
  assign _0566_ = _0507_ & _0104_;
  assign _0564_ = _0508_ & _0104_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) md_state_q <= 3'h0;
    else if (div_en_internal) md_state_q <= md_state_d;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) div_counter_q <= 5'h00;
    else if (div_en_internal) div_counter_q <= div_counter_d;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) \gen_mult_single_cycle.mult_state_q  <= 1'h0;
    else if (mult_en_internal) \gen_mult_single_cycle.mult_state_q  <= \gen_mult_single_cycle.mult_state_d ;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) op_quotient_q <= 32'd0;
    else if (_0020_) op_quotient_q <= op_quotient_d;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) op_numerator_q <= 32'd0;
    else if (_0022_) op_numerator_q <= _0573_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) div_by_zero_q <= 1'h0;
    else if (_0024_) div_by_zero_q <= equal_to_zero_i;
  assign _0227_ = data_ind_timing_i_t0 & equal_to_zero_i;
  assign _0228_ = equal_to_zero_i_t0 & _0546_;
  assign _0229_ = data_ind_timing_i_t0 & equal_to_zero_i_t0;
  assign _0403_ = _0227_ | _0228_;
  assign _0545_ = _0403_ | _0229_;
  assign _0094_ = | { _0568_, _0566_ };
  assign _0098_ = | { _0560_, _0568_ };
  assign _0099_ = | { _0564_, _0562_, _0566_ };
  assign _0100_ = | { _0558_, _0560_, _0568_ };
  assign _0103_ = | signed_mode_i_t0;
  assign _0102_ = | operator_i_t0;
  assign _0038_ = ~ { _0568_, _0566_ };
  assign _0039_ = ~ { _0568_, _0560_ };
  assign _0040_ = ~ { _0566_, _0564_, _0562_ };
  assign _0045_ = ~ { _0568_, _0560_, _0558_ };
  assign _0065_ = ~ signed_mode_i_t0;
  assign _0153_ = { _0567_, _0565_ } & _0038_;
  assign _0154_ = { _0567_, _0559_ } & _0039_;
  assign _0155_ = { _0565_, _0563_, _0561_ } & _0040_;
  assign _0162_ = { _0567_, _0559_, _0557_ } & _0045_;
  assign _0230_ = signed_mode_i & _0065_;
  assign _0106_ = ! _0153_;
  assign _0107_ = ! _0154_;
  assign _0108_ = ! _0155_;
  assign _0109_ = ! _0162_;
  assign _0110_ = ! _0230_;
  assign _0111_ = ! _0225_;
  assign _0112_ = ! _0262_;
  assign _0019_ = _0106_ & _0094_;
  assign _0027_ = _0107_ & _0098_;
  assign _0029_ = _0108_ & _0099_;
  assign _0093_ = _0109_ & _0100_;
  assign signed_mult_t0 = _0110_ & _0103_;
  assign _0001_ = _0111_ & _0102_;
  assign _0562_ = _0112_ & _0104_;
  assign _0047_ = ~ { \gen_mult_single_cycle.mult_state_q , \gen_mult_single_cycle.mult_state_q , \gen_mult_single_cycle.mult_state_q , \gen_mult_single_cycle.mult_state_q , \gen_mult_single_cycle.mult_state_q , \gen_mult_single_cycle.mult_state_q , \gen_mult_single_cycle.mult_state_q , \gen_mult_single_cycle.mult_state_q , \gen_mult_single_cycle.mult_state_q , \gen_mult_single_cycle.mult_state_q , \gen_mult_single_cycle.mult_state_q , \gen_mult_single_cycle.mult_state_q , \gen_mult_single_cycle.mult_state_q , \gen_mult_single_cycle.mult_state_q , \gen_mult_single_cycle.mult_state_q , \gen_mult_single_cycle.mult_state_q , \gen_mult_single_cycle.mult_state_q , \gen_mult_single_cycle.mult_state_q , \gen_mult_single_cycle.mult_state_q , \gen_mult_single_cycle.mult_state_q , \gen_mult_single_cycle.mult_state_q , \gen_mult_single_cycle.mult_state_q , \gen_mult_single_cycle.mult_state_q , \gen_mult_single_cycle.mult_state_q , \gen_mult_single_cycle.mult_state_q , \gen_mult_single_cycle.mult_state_q , \gen_mult_single_cycle.mult_state_q , \gen_mult_single_cycle.mult_state_q , \gen_mult_single_cycle.mult_state_q , \gen_mult_single_cycle.mult_state_q , \gen_mult_single_cycle.mult_state_q , \gen_mult_single_cycle.mult_state_q , \gen_mult_single_cycle.mult_state_q , \gen_mult_single_cycle.mult_state_q  };
  assign _0046_ = ~ \gen_mult_single_cycle.mult_state_q ;
  assign _0048_ = ~ { _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_ };
  assign _0049_ = ~ { _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_ };
  assign _0050_ = ~ { _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_ };
  assign _0051_ = ~ { _0559_, _0559_, _0559_ };
  assign _0052_ = ~ { _0557_, _0557_, _0557_ };
  assign _0053_ = ~ { _0563_, _0563_, _0563_ };
  assign _0054_ = ~ { _0561_, _0561_, _0561_ };
  assign _0055_ = ~ { _0309_, _0309_, _0309_ };
  assign _0056_ = ~ { _0092_, _0092_, _0092_ };
  assign _0057_ = ~ { _0559_, _0559_, _0559_, _0559_, _0559_, _0559_, _0559_, _0559_, _0559_, _0559_, _0559_, _0559_, _0559_, _0559_, _0559_, _0559_, _0559_, _0559_, _0559_, _0559_, _0559_, _0559_, _0559_, _0559_, _0559_, _0559_, _0559_, _0559_, _0559_, _0559_, _0559_, _0559_, _0559_, _0559_ };
  assign _0058_ = ~ { _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_ };
  assign _0059_ = ~ { _0561_, _0561_, _0561_, _0561_, _0561_, _0561_, _0561_, _0561_, _0561_, _0561_, _0561_, _0561_, _0561_, _0561_, _0561_, _0561_, _0561_, _0561_, _0561_, _0561_, _0561_, _0561_, _0561_, _0561_, _0561_, _0561_, _0561_, _0561_, _0561_, _0561_, _0561_, _0561_, _0561_, _0561_ };
  assign _0060_ = ~ { _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_ };
  assign _0061_ = ~ { _0092_, _0092_, _0092_, _0092_, _0092_, _0092_, _0092_, _0092_, _0092_, _0092_, _0092_, _0092_, _0092_, _0092_, _0092_, _0092_, _0092_, _0092_, _0092_, _0092_, _0092_, _0092_, _0092_, _0092_, _0092_, _0092_, _0092_, _0092_, _0092_, _0092_, _0092_, _0092_, _0092_, _0092_ };
  assign _0062_ = ~ { _0567_, _0567_, _0567_, _0567_, _0567_, _0567_, _0567_, _0567_, _0567_, _0567_, _0567_, _0567_, _0567_, _0567_, _0567_, _0567_, _0567_, _0567_, _0567_, _0567_, _0567_, _0567_, _0567_, _0567_, _0567_, _0567_, _0567_, _0567_, _0567_, _0567_, _0567_, _0567_ };
  assign _0071_ = ~ { _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_ };
  assign _0070_ = ~ _0547_;
  assign _0072_ = ~ { _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_ };
  assign _0073_ = ~ { _0028_, _0028_, _0028_, _0028_, _0028_ };
  assign _0074_ = ~ { _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_ };
  assign _0076_ = ~ { _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_ };
  assign _0077_ = ~ _0583_;
  assign _0078_ = ~ { div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i };
  assign _0079_ = ~ { div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i };
  assign _0080_ = ~ { is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal };
  assign _0081_ = ~ { is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal };
  assign _0082_ = ~ { _0544_, _0544_, _0544_ };
  assign _0083_ = ~ { div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a };
  assign _0084_ = ~ { div_sign_b, div_sign_b, div_sign_b, div_sign_b, div_sign_b, div_sign_b, div_sign_b, div_sign_b, div_sign_b, div_sign_b, div_sign_b, div_sign_b, div_sign_b, div_sign_b, div_sign_b, div_sign_b, div_sign_b, div_sign_b, div_sign_b, div_sign_b, div_sign_b, div_sign_b, div_sign_b, div_sign_b, div_sign_b, div_sign_b, div_sign_b, div_sign_b, div_sign_b, div_sign_b, div_sign_b, div_sign_b };
  assign _0085_ = ~ { _0542_, _0542_, _0542_ };
  assign _0086_ = ~ { div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign };
  assign _0087_ = ~ { div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a };
  assign _0353_ = { \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0  } | _0047_;
  assign _0350_ = \gen_mult_single_cycle.mult_state_q_t0  | _0046_;
  assign _0358_ = { _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_ } | _0048_;
  assign _0361_ = { _0566_, _0566_, _0566_, _0566_, _0566_, _0566_, _0566_, _0566_, _0566_, _0566_, _0566_, _0566_, _0566_, _0566_, _0566_, _0566_, _0566_, _0566_, _0566_, _0566_, _0566_, _0566_, _0566_, _0566_, _0566_, _0566_, _0566_, _0566_, _0566_, _0566_, _0566_, _0566_, _0566_ } | _0049_;
  assign _0364_ = { _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_ } | _0050_;
  assign _0367_ = { _0560_, _0560_, _0560_ } | _0051_;
  assign _0370_ = { _0558_, _0558_, _0558_ } | _0052_;
  assign _0373_ = { _0564_, _0564_, _0564_ } | _0053_;
  assign _0376_ = { _0562_, _0562_, _0562_ } | _0054_;
  assign _0379_ = { _0310_, _0310_, _0310_ } | _0055_;
  assign _0382_ = { _0093_, _0093_, _0093_ } | _0056_;
  assign _0385_ = { _0560_, _0560_, _0560_, _0560_, _0560_, _0560_, _0560_, _0560_, _0560_, _0560_, _0560_, _0560_, _0560_, _0560_, _0560_, _0560_, _0560_, _0560_, _0560_, _0560_, _0560_, _0560_, _0560_, _0560_, _0560_, _0560_, _0560_, _0560_, _0560_, _0560_, _0560_, _0560_, _0560_, _0560_ } | _0057_;
  assign _0388_ = { _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_ } | _0058_;
  assign _0391_ = { _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_ } | _0059_;
  assign _0394_ = { _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_ } | _0060_;
  assign _0397_ = { _0093_, _0093_, _0093_, _0093_, _0093_, _0093_, _0093_, _0093_, _0093_, _0093_, _0093_, _0093_, _0093_, _0093_, _0093_, _0093_, _0093_, _0093_, _0093_, _0093_, _0093_, _0093_, _0093_, _0093_, _0093_, _0093_, _0093_, _0093_, _0093_, _0093_, _0093_, _0093_, _0093_, _0093_ } | _0061_;
  assign _0400_ = { _0568_, _0568_, _0568_, _0568_, _0568_, _0568_, _0568_, _0568_, _0568_, _0568_, _0568_, _0568_, _0568_, _0568_, _0568_, _0568_, _0568_, _0568_, _0568_, _0568_, _0568_, _0568_, _0568_, _0568_, _0568_, _0568_, _0568_, _0568_, _0568_, _0568_, _0568_, _0568_ } | _0062_;
  assign _0408_ = { _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_ } | _0071_;
  assign _0407_ = _0001_ | _0070_;
  assign _0411_ = { _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_ } | _0072_;
  assign _0416_ = { _0029_, _0029_, _0029_, _0029_, _0029_ } | _0073_;
  assign _0419_ = { _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_ } | _0074_;
  assign _0423_ = { _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_ } | _0076_;
  assign _0426_ = _0584_ | _0077_;
  assign _0431_ = { div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0 } | _0078_;
  assign _0434_ = { div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0 } | _0079_;
  assign _0437_ = { is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0 } | _0080_;
  assign _0440_ = { is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0 } | _0081_;
  assign _0443_ = { _0545_, _0545_, _0545_ } | _0082_;
  assign _0446_ = { div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0 } | _0083_;
  assign _0449_ = { div_sign_b_t0, div_sign_b_t0, div_sign_b_t0, div_sign_b_t0, div_sign_b_t0, div_sign_b_t0, div_sign_b_t0, div_sign_b_t0, div_sign_b_t0, div_sign_b_t0, div_sign_b_t0, div_sign_b_t0, div_sign_b_t0, div_sign_b_t0, div_sign_b_t0, div_sign_b_t0, div_sign_b_t0, div_sign_b_t0, div_sign_b_t0, div_sign_b_t0, div_sign_b_t0, div_sign_b_t0, div_sign_b_t0, div_sign_b_t0, div_sign_b_t0, div_sign_b_t0, div_sign_b_t0, div_sign_b_t0, div_sign_b_t0, div_sign_b_t0, div_sign_b_t0, div_sign_b_t0 } | _0084_;
  assign _0452_ = { _0543_, _0543_, _0543_ } | _0085_;
  assign _0455_ = { div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0 } | _0086_;
  assign _0458_ = { div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0 } | _0087_;
  assign _0354_ = { \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0  } | { \gen_mult_single_cycle.mult_state_q , \gen_mult_single_cycle.mult_state_q , \gen_mult_single_cycle.mult_state_q , \gen_mult_single_cycle.mult_state_q , \gen_mult_single_cycle.mult_state_q , \gen_mult_single_cycle.mult_state_q , \gen_mult_single_cycle.mult_state_q , \gen_mult_single_cycle.mult_state_q , \gen_mult_single_cycle.mult_state_q , \gen_mult_single_cycle.mult_state_q , \gen_mult_single_cycle.mult_state_q , \gen_mult_single_cycle.mult_state_q , \gen_mult_single_cycle.mult_state_q , \gen_mult_single_cycle.mult_state_q , \gen_mult_single_cycle.mult_state_q , \gen_mult_single_cycle.mult_state_q , \gen_mult_single_cycle.mult_state_q , \gen_mult_single_cycle.mult_state_q , \gen_mult_single_cycle.mult_state_q , \gen_mult_single_cycle.mult_state_q , \gen_mult_single_cycle.mult_state_q , \gen_mult_single_cycle.mult_state_q , \gen_mult_single_cycle.mult_state_q , \gen_mult_single_cycle.mult_state_q , \gen_mult_single_cycle.mult_state_q , \gen_mult_single_cycle.mult_state_q , \gen_mult_single_cycle.mult_state_q , \gen_mult_single_cycle.mult_state_q , \gen_mult_single_cycle.mult_state_q , \gen_mult_single_cycle.mult_state_q , \gen_mult_single_cycle.mult_state_q , \gen_mult_single_cycle.mult_state_q , \gen_mult_single_cycle.mult_state_q , \gen_mult_single_cycle.mult_state_q  };
  assign _0351_ = \gen_mult_single_cycle.mult_state_q_t0  | \gen_mult_single_cycle.mult_state_q ;
  assign _0359_ = { _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_ } | { _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_ };
  assign _0362_ = { _0566_, _0566_, _0566_, _0566_, _0566_, _0566_, _0566_, _0566_, _0566_, _0566_, _0566_, _0566_, _0566_, _0566_, _0566_, _0566_, _0566_, _0566_, _0566_, _0566_, _0566_, _0566_, _0566_, _0566_, _0566_, _0566_, _0566_, _0566_, _0566_, _0566_, _0566_, _0566_, _0566_ } | { _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_ };
  assign _0365_ = { _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_ } | { _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_ };
  assign _0368_ = { _0560_, _0560_, _0560_ } | { _0559_, _0559_, _0559_ };
  assign _0371_ = { _0558_, _0558_, _0558_ } | { _0557_, _0557_, _0557_ };
  assign _0374_ = { _0564_, _0564_, _0564_ } | { _0563_, _0563_, _0563_ };
  assign _0377_ = { _0562_, _0562_, _0562_ } | { _0561_, _0561_, _0561_ };
  assign _0380_ = { _0310_, _0310_, _0310_ } | { _0309_, _0309_, _0309_ };
  assign _0383_ = { _0093_, _0093_, _0093_ } | { _0092_, _0092_, _0092_ };
  assign _0386_ = { _0560_, _0560_, _0560_, _0560_, _0560_, _0560_, _0560_, _0560_, _0560_, _0560_, _0560_, _0560_, _0560_, _0560_, _0560_, _0560_, _0560_, _0560_, _0560_, _0560_, _0560_, _0560_, _0560_, _0560_, _0560_, _0560_, _0560_, _0560_, _0560_, _0560_, _0560_, _0560_, _0560_, _0560_ } | { _0559_, _0559_, _0559_, _0559_, _0559_, _0559_, _0559_, _0559_, _0559_, _0559_, _0559_, _0559_, _0559_, _0559_, _0559_, _0559_, _0559_, _0559_, _0559_, _0559_, _0559_, _0559_, _0559_, _0559_, _0559_, _0559_, _0559_, _0559_, _0559_, _0559_, _0559_, _0559_, _0559_, _0559_ };
  assign _0389_ = { _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_ } | { _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_ };
  assign _0392_ = { _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_ } | { _0561_, _0561_, _0561_, _0561_, _0561_, _0561_, _0561_, _0561_, _0561_, _0561_, _0561_, _0561_, _0561_, _0561_, _0561_, _0561_, _0561_, _0561_, _0561_, _0561_, _0561_, _0561_, _0561_, _0561_, _0561_, _0561_, _0561_, _0561_, _0561_, _0561_, _0561_, _0561_, _0561_, _0561_ };
  assign _0395_ = { _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_ } | { _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_ };
  assign _0398_ = { _0093_, _0093_, _0093_, _0093_, _0093_, _0093_, _0093_, _0093_, _0093_, _0093_, _0093_, _0093_, _0093_, _0093_, _0093_, _0093_, _0093_, _0093_, _0093_, _0093_, _0093_, _0093_, _0093_, _0093_, _0093_, _0093_, _0093_, _0093_, _0093_, _0093_, _0093_, _0093_, _0093_, _0093_ } | { _0092_, _0092_, _0092_, _0092_, _0092_, _0092_, _0092_, _0092_, _0092_, _0092_, _0092_, _0092_, _0092_, _0092_, _0092_, _0092_, _0092_, _0092_, _0092_, _0092_, _0092_, _0092_, _0092_, _0092_, _0092_, _0092_, _0092_, _0092_, _0092_, _0092_, _0092_, _0092_, _0092_, _0092_ };
  assign _0401_ = { _0568_, _0568_, _0568_, _0568_, _0568_, _0568_, _0568_, _0568_, _0568_, _0568_, _0568_, _0568_, _0568_, _0568_, _0568_, _0568_, _0568_, _0568_, _0568_, _0568_, _0568_, _0568_, _0568_, _0568_, _0568_, _0568_, _0568_, _0568_, _0568_, _0568_, _0568_, _0568_ } | { _0567_, _0567_, _0567_, _0567_, _0567_, _0567_, _0567_, _0567_, _0567_, _0567_, _0567_, _0567_, _0567_, _0567_, _0567_, _0567_, _0567_, _0567_, _0567_, _0567_, _0567_, _0567_, _0567_, _0567_, _0567_, _0567_, _0567_, _0567_, _0567_, _0567_, _0567_, _0567_ };
  assign _0409_ = { _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_ } | { _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_ };
  assign _0412_ = { _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_ } | { _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_ };
  assign _0417_ = { _0029_, _0029_, _0029_, _0029_, _0029_ } | { _0028_, _0028_, _0028_, _0028_, _0028_ };
  assign _0420_ = { _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_ } | { _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_ };
  assign _0422_ = div_valid_t0 | _0569_;
  assign _0424_ = { _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_ } | { _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_ };
  assign _0427_ = _0584_ | _0583_;
  assign _0432_ = { div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0 } | { div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i };
  assign _0435_ = { div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0 } | { div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i, div_sel_i };
  assign _0438_ = { is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0 } | { is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal };
  assign _0441_ = { is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0 } | { is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal };
  assign _0444_ = { _0545_, _0545_, _0545_ } | { _0544_, _0544_, _0544_ };
  assign _0447_ = { div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0 } | { div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a };
  assign _0450_ = { div_sign_b_t0, div_sign_b_t0, div_sign_b_t0, div_sign_b_t0, div_sign_b_t0, div_sign_b_t0, div_sign_b_t0, div_sign_b_t0, div_sign_b_t0, div_sign_b_t0, div_sign_b_t0, div_sign_b_t0, div_sign_b_t0, div_sign_b_t0, div_sign_b_t0, div_sign_b_t0, div_sign_b_t0, div_sign_b_t0, div_sign_b_t0, div_sign_b_t0, div_sign_b_t0, div_sign_b_t0, div_sign_b_t0, div_sign_b_t0, div_sign_b_t0, div_sign_b_t0, div_sign_b_t0, div_sign_b_t0, div_sign_b_t0, div_sign_b_t0, div_sign_b_t0, div_sign_b_t0 } | { div_sign_b, div_sign_b, div_sign_b, div_sign_b, div_sign_b, div_sign_b, div_sign_b, div_sign_b, div_sign_b, div_sign_b, div_sign_b, div_sign_b, div_sign_b, div_sign_b, div_sign_b, div_sign_b, div_sign_b, div_sign_b, div_sign_b, div_sign_b, div_sign_b, div_sign_b, div_sign_b, div_sign_b, div_sign_b, div_sign_b, div_sign_b, div_sign_b, div_sign_b, div_sign_b, div_sign_b, div_sign_b };
  assign _0453_ = { _0543_, _0543_, _0543_ } | { _0542_, _0542_, _0542_ };
  assign _0456_ = { div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0 } | { div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign };
  assign _0459_ = { div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0 } | { div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a };
  assign _0163_ = _0001_ & _0350_;
  assign _0165_ = _0007_ & _0350_;
  assign _0168_ = _0003_ & _0353_;
  assign _0171_ = _0009_ & _0350_;
  assign _0173_ = 34'h000000000 & _0353_;
  assign _0178_ = { imd_val_q_i_t0[31:0], 1'h0 } & _0358_;
  assign _0181_ = { op_b_i_t0, 1'h0 } & _0361_;
  assign _0184_ = _0518_ & _0364_;
  assign _0187_ = _0578_ & _0367_;
  assign _0190_ = _0520_ & _0370_;
  assign _0193_ = 3'h0 & _0373_;
  assign _0196_ = 3'h0 & _0376_;
  assign _0199_ = _0526_ & _0379_;
  assign _0202_ = _0528_ & _0382_;
  assign _0205_ = { 1'h0, next_remainder_t0, _0571_ } & _0385_;
  assign _0208_ = _0530_ & _0388_;
  assign _0211_ = imd_val_q_i_t0[67:34] & _0391_;
  assign _0214_ = _0534_ & _0394_;
  assign _0217_ = _0536_ & _0397_;
  assign _0220_ = 32'd0 & _0400_;
  assign _0240_ = mult_en_i_t0 & _0407_;
  assign _0242_ = { 2'h0, mac_res_ext_t0[15:0], 16'h0000 } & _0408_;
  assign _0245_ = multdiv_ready_id_i_t0 & _0407_;
  assign _0247_ = _0582_ & _0411_;
  assign _0250_ = { 2'h0, next_remainder_t0 } & _0411_;
  assign _0253_ = { 2'h0, op_a_i_t0 } & _0411_;
  assign _0256_ = _0430_ & _0416_;
  assign _0259_ = 33'h000000000 & _0419_;
  assign _0270_ = imd_val_q_i_t0[31:0] & _0423_;
  assign _0274_ = alu_adder_ext_i_t0[32] & _0426_;
  assign _0277_ = mac_res_d_t0 & _0431_;
  assign _0280_ = mac_res_d_t0[31:0] & _0434_;
  assign _0283_ = imd_val_q_i_t0[65:34] & _0437_;
  assign _0286_ = { 1'h0, op_quotient_q_t0 } & _0440_;
  assign _0289_ = 3'h0 & _0443_;
  assign _0292_ = op_a_i_t0 & _0446_;
  assign _0295_ = op_b_i_t0 & _0449_;
  assign _0298_ = 3'h0 & _0452_;
  assign _0301_ = imd_val_q_i_t0[67:34] & _0455_;
  assign _0304_ = imd_val_q_i_t0[67:34] & _0458_;
  assign _0166_ = multdiv_ready_id_i_t0 & _0351_;
  assign _0169_ = mac_res_ext_t0[33:0] & _0354_;
  assign _0174_ = { accum_t0[33], accum_t0[33], accum_t0[33], accum_t0[33], accum_t0[33], accum_t0[33], accum_t0[33], accum_t0[33], accum_t0[33], accum_t0[33], accum_t0[33], accum_t0[33], accum_t0[33], accum_t0[33], accum_t0[33], accum_t0[33], imd_val_q_i_t0[67:50] } & _0354_;
  assign _0176_ = 34'h000000000 & _0354_;
  assign _0179_ = { imd_val_q_i_t0[65:34], 1'h0 } & _0359_;
  assign _0182_ = { op_a_i_t0, 1'h0 } & _0362_;
  assign _0185_ = _0516_ & _0365_;
  assign _0188_ = 3'h0 & _0368_;
  assign _0191_ = 3'h0 & _0371_;
  assign _0194_ = 3'h0 & _0374_;
  assign _0197_ = _0005_ & _0377_;
  assign _0200_ = _0524_ & _0380_;
  assign _0203_ = _0522_ & _0383_;
  assign _0206_ = _0013_ & _0386_;
  assign _0209_ = _0015_ & _0389_;
  assign _0212_ = _0011_ & _0392_;
  assign _0215_ = { 33'h000000000, op_numerator_q_t0[31] } & _0395_;
  assign _0218_ = _0532_ & _0398_;
  assign _0221_ = next_quotient_t0[31:0] & _0401_;
  assign _0243_ = mac_res_ext_t0[33:0] & _0409_;
  assign _0248_ = _0580_ & _0412_;
  assign _0251_ = { 1'h0, next_quotient_t0 } & _0412_;
  assign _0254_ = 34'h000000000 & _0412_;
  assign _0257_ = 5'h00 & _0417_;
  assign _0260_ = { imd_val_q_i_t0[65:34], 1'h0 } & _0420_;
  assign _0265_ = multdiv_ready_id_i_t0 & _0422_;
  assign _0271_ = _0576_ & _0424_;
  assign _0275_ = imd_val_q_i_t0[65] & _0427_;
  assign _0278_ = op_remainder_d_t0 & _0432_;
  assign _0281_ = imd_val_q_i_t0[65:34] & _0435_;
  assign _0284_ = alu_adder_ext_i_t0[32:1] & _0438_;
  assign _0287_ = _0556_ & _0441_;
  assign _0290_ = 3'h0 & _0444_;
  assign _0293_ = alu_adder_i_t0 & _0447_;
  assign _0296_ = alu_adder_i_t0 & _0450_;
  assign _0299_ = 3'h0 & _0453_;
  assign _0302_ = { 2'h0, alu_adder_i_t0 } & _0456_;
  assign _0305_ = { 2'h0, alu_adder_i_t0 } & _0459_;
  assign _0352_ = _0165_ | _0166_;
  assign _0355_ = _0168_ | _0169_;
  assign _0356_ = _0173_ | _0174_;
  assign _0357_ = _0173_ | _0176_;
  assign _0360_ = _0178_ | _0179_;
  assign _0363_ = _0181_ | _0182_;
  assign _0366_ = _0184_ | _0185_;
  assign _0369_ = _0187_ | _0188_;
  assign _0372_ = _0190_ | _0191_;
  assign _0375_ = _0193_ | _0194_;
  assign _0378_ = _0196_ | _0197_;
  assign _0381_ = _0199_ | _0200_;
  assign _0384_ = _0202_ | _0203_;
  assign _0387_ = _0205_ | _0206_;
  assign _0390_ = _0208_ | _0209_;
  assign _0393_ = _0211_ | _0212_;
  assign _0396_ = _0214_ | _0215_;
  assign _0399_ = _0217_ | _0218_;
  assign _0402_ = _0220_ | _0221_;
  assign _0410_ = _0242_ | _0243_;
  assign _0413_ = _0247_ | _0248_;
  assign _0414_ = _0250_ | _0251_;
  assign _0415_ = _0253_ | _0254_;
  assign _0418_ = _0256_ | _0257_;
  assign _0421_ = _0259_ | _0260_;
  assign _0425_ = _0270_ | _0271_;
  assign _0428_ = _0274_ | _0275_;
  assign _0433_ = _0277_ | _0278_;
  assign _0436_ = _0280_ | _0281_;
  assign _0439_ = _0283_ | _0284_;
  assign _0442_ = _0286_ | _0287_;
  assign _0445_ = _0289_ | _0290_;
  assign _0448_ = _0292_ | _0293_;
  assign _0451_ = _0295_ | _0296_;
  assign _0454_ = _0298_ | _0299_;
  assign _0457_ = _0301_ | _0302_;
  assign _0460_ = _0304_ | _0305_;
  assign _0469_ = _0006_ ^ _0485_;
  assign _0470_ = _0002_ ^ mac_res_ext[33:0];
  assign _0471_ = \gen_mult_single_cycle.mult2_res  ^ { accum[33], accum[33], accum[33], accum[33], accum[33], accum[33], accum[33], accum[33], accum[33], accum[33], accum[33], accum[33], accum[33], accum[33], accum[33], accum[33], imd_val_q_i[67:50] };
  assign _0472_ = { _0553_, 1'h1 } ^ { _0554_, 1'h1 };
  assign _0473_ = { _0551_, 1'h1 } ^ { _0552_, 1'h1 };
  assign _0474_ = _0517_ ^ _0515_;
  assign _0475_ = _0577_ ^ 3'h5;
  assign _0476_ = _0519_ ^ 3'h6;
  assign _0477_ = _0525_ ^ _0523_;
  assign _0478_ = _0527_ ^ _0521_;
  assign _0479_ = { 1'h0, next_remainder, _0570_ } ^ _0012_;
  assign _0480_ = _0529_ ^ _0014_;
  assign _0481_ = imd_val_q_i[67:34] ^ _0010_;
  assign _0482_ = _0533_ ^ { 33'h000000000, op_numerator_q[31] };
  assign _0483_ = _0535_ ^ _0531_;
  assign _0484_ = { 2'h0, mac_res_ext[15:0], \gen_mult_single_cycle.mult1_res [15:0] } ^ mac_res_ext[33:0];
  assign _0486_ = _0581_ ^ _0579_;
  assign _0487_ = { 2'h0, next_remainder } ^ { 1'h0, next_quotient };
  assign _0488_ = { 2'h0, op_a_i } ^ 34'h3ffffffff;
  assign _0489_ = _0572_ ^ 5'h1f;
  assign _0490_ = 33'h000000001 ^ { imd_val_q_i[65:34], 1'h1 };
  assign _0491_ = imd_val_q_i[31:0] ^ _0575_;
  assign _0492_ = _0539_ ^ imd_val_q_i[65];
  assign _0494_ = mac_res_d ^ op_remainder_d;
  assign _0495_ = mac_res_d[31:0] ^ imd_val_q_i[65:34];
  assign _0496_ = imd_val_q_i[65:34] ^ alu_adder_ext_i[32:1];
  assign _0497_ = { 1'h0, op_quotient_q } ^ _0555_;
  assign _0498_ = op_a_i ^ alu_adder_i;
  assign _0499_ = op_b_i ^ alu_adder_i;
  assign _0500_ = imd_val_q_i[67:34] ^ { 2'h0, alu_adder_i };
  assign _0164_ = \gen_mult_single_cycle.mult_state_q_t0  & _0000_;
  assign _0167_ = \gen_mult_single_cycle.mult_state_q_t0  & _0469_;
  assign _0170_ = { \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0  } & _0470_;
  assign _0172_ = \gen_mult_single_cycle.mult_state_q_t0  & _0088_;
  assign _0175_ = { \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0  } & _0471_;
  assign _0177_ = { \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0 , \gen_mult_single_cycle.mult_state_q_t0  } & { 18'h00000, \gen_mult_single_cycle.mult1_res [31:16] };
  assign _0180_ = { _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_ } & _0472_;
  assign _0183_ = { _0566_, _0566_, _0566_, _0566_, _0566_, _0566_, _0566_, _0566_, _0566_, _0566_, _0566_, _0566_, _0566_, _0566_, _0566_, _0566_, _0566_, _0566_, _0566_, _0566_, _0566_, _0566_, _0566_, _0566_, _0566_, _0566_, _0566_, _0566_, _0566_, _0566_, _0566_, _0566_, _0566_ } & _0473_;
  assign _0186_ = { _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_ } & _0474_;
  assign _0189_ = { _0560_, _0560_, _0560_ } & _0475_;
  assign _0192_ = { _0558_, _0558_, _0558_ } & _0476_;
  assign _0195_ = { _0564_, _0564_, _0564_ } & 3'h1;
  assign _0198_ = { _0562_, _0562_, _0562_ } & _0004_;
  assign _0201_ = { _0310_, _0310_, _0310_ } & _0477_;
  assign _0204_ = { _0093_, _0093_, _0093_ } & _0478_;
  assign _0207_ = { _0560_, _0560_, _0560_, _0560_, _0560_, _0560_, _0560_, _0560_, _0560_, _0560_, _0560_, _0560_, _0560_, _0560_, _0560_, _0560_, _0560_, _0560_, _0560_, _0560_, _0560_, _0560_, _0560_, _0560_, _0560_, _0560_, _0560_, _0560_, _0560_, _0560_, _0560_, _0560_, _0560_, _0560_ } & _0479_;
  assign _0210_ = { _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_, _0558_ } & _0480_;
  assign _0213_ = { _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_ } & _0481_;
  assign _0216_ = { _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_ } & _0482_;
  assign _0219_ = { _0093_, _0093_, _0093_, _0093_, _0093_, _0093_, _0093_, _0093_, _0093_, _0093_, _0093_, _0093_, _0093_, _0093_, _0093_, _0093_, _0093_, _0093_, _0093_, _0093_, _0093_, _0093_, _0093_, _0093_, _0093_, _0093_, _0093_, _0093_, _0093_, _0093_, _0093_, _0093_, _0093_, _0093_ } & _0483_;
  assign _0222_ = { _0568_, _0568_, _0568_, _0568_, _0568_, _0568_, _0568_, _0568_, _0568_, _0568_, _0568_, _0568_, _0568_, _0568_, _0568_, _0568_, _0568_, _0568_, _0568_, _0568_, _0568_, _0568_, _0568_, _0568_, _0568_, _0568_, _0568_, _0568_, _0568_, _0568_, _0568_, _0568_ } & next_quotient[31:0];
  assign _0241_ = _0001_ & mult_en_i;
  assign _0244_ = { _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_ } & _0484_;
  assign _0246_ = _0001_ & _0485_;
  assign _0249_ = { _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_ } & _0486_;
  assign _0252_ = { _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_ } & _0487_;
  assign _0255_ = { _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_ } & _0488_;
  assign _0258_ = { _0029_, _0029_, _0029_, _0029_, _0029_ } & _0489_;
  assign _0261_ = { _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_ } & _0490_;
  assign _0266_ = div_valid_t0 & _0485_;
  assign _0272_ = { _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_ } & _0491_;
  assign _0276_ = _0584_ & _0492_;
  assign _0279_ = { div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0 } & _0494_;
  assign _0282_ = { div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0, div_sel_i_t0 } & _0495_;
  assign _0285_ = { is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0 } & _0496_;
  assign _0288_ = { is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0 } & _0497_;
  assign _0291_ = { _0545_, _0545_, _0545_ } & 3'h7;
  assign _0294_ = { div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0 } & _0498_;
  assign _0297_ = { div_sign_b_t0, div_sign_b_t0, div_sign_b_t0, div_sign_b_t0, div_sign_b_t0, div_sign_b_t0, div_sign_b_t0, div_sign_b_t0, div_sign_b_t0, div_sign_b_t0, div_sign_b_t0, div_sign_b_t0, div_sign_b_t0, div_sign_b_t0, div_sign_b_t0, div_sign_b_t0, div_sign_b_t0, div_sign_b_t0, div_sign_b_t0, div_sign_b_t0, div_sign_b_t0, div_sign_b_t0, div_sign_b_t0, div_sign_b_t0, div_sign_b_t0, div_sign_b_t0, div_sign_b_t0, div_sign_b_t0, div_sign_b_t0, div_sign_b_t0, div_sign_b_t0, div_sign_b_t0 } & _0499_;
  assign _0300_ = { _0543_, _0543_, _0543_ } & 3'h7;
  assign _0303_ = { div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0 } & _0500_;
  assign _0306_ = { div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0, div_sign_a_t0 } & _0500_;
  assign \gen_mult_single_cycle.mult_state_d_t0  = _0164_ | _0163_;
  assign mult_hold_t0 = _0167_ | _0352_;
  assign mac_res_d_t0 = _0170_ | _0355_;
  assign mult_valid_t0 = _0172_ | _0171_;
  assign \gen_mult_single_cycle.summand2_t0  = _0175_ | _0356_;
  assign \gen_mult_single_cycle.summand1_t0  = _0177_ | _0357_;
  assign _0516_ = _0180_ | _0360_;
  assign _0518_ = _0183_ | _0363_;
  assign alu_operand_b_o_t0 = _0186_ | _0366_;
  assign _0520_ = _0189_ | _0369_;
  assign _0522_ = _0192_ | _0372_;
  assign _0524_ = _0195_ | _0375_;
  assign _0526_ = _0198_ | _0378_;
  assign _0528_ = _0201_ | _0381_;
  assign md_state_d_t0 = _0204_ | _0384_;
  assign _0530_ = _0207_ | _0387_;
  assign _0532_ = _0210_ | _0390_;
  assign _0534_ = _0213_ | _0393_;
  assign _0536_ = _0216_ | _0396_;
  assign op_remainder_d_t0 = _0219_ | _0399_;
  assign op_quotient_d_t0 = _0222_ | _0402_;
  assign _0009_ = _0241_ | _0240_;
  assign _0003_ = _0244_ | _0410_;
  assign _0007_ = _0246_ | _0245_;
  assign _0015_ = _0249_ | _0413_;
  assign _0013_ = _0252_ | _0414_;
  assign _0011_ = _0255_ | _0415_;
  assign div_counter_d_t0 = _0258_ | _0418_;
  assign alu_operand_a_o_t0 = _0261_ | _0421_;
  assign div_hold_t0 = _0266_ | _0265_;
  assign op_denominator_d_t0 = _0272_ | _0425_;
  assign is_greater_equal_t0 = _0276_ | _0428_;
  assign imd_val_d_o_t0[67:34] = _0279_ | _0433_;
  assign multdiv_result_o_t0 = _0282_ | _0436_;
  assign next_remainder_t0 = _0285_ | _0439_;
  assign next_quotient_t0 = _0288_ | _0442_;
  assign _0005_ = _0291_ | _0445_;
  assign _0574_ = _0294_ | _0448_;
  assign _0576_ = _0297_ | _0451_;
  assign _0578_ = _0300_ | _0454_;
  assign _0580_ = _0303_ | _0457_;
  assign _0582_ = _0306_ | _0460_;
  assign _0018_ = | { _0567_, _0565_ };
  assign _0020_ = & { _0018_, div_en_internal };
  assign _0022_ = & { _0565_, div_en_internal };
  assign _0024_ = & { _0561_, _0540_, div_en_internal };
  assign _0088_ = ~ _0008_;
  assign _0026_ = | { _0567_, _0559_ };
  assign _0028_ = | { _0565_, _0563_, _0561_ };
  assign _0041_ = ~ _0026_;
  assign _0043_ = ~ _0565_;
  assign _0034_ = ~ mult_en_internal;
  assign _0066_ = ~ { 1'h0, op_quotient_q };
  assign _0068_ = ~ mult_valid;
  assign _0042_ = ~ _0557_;
  assign _0044_ = ~ _0563_;
  assign _0033_ = ~ div_en_internal;
  assign _0067_ = ~ { 1'h0, one_shift };
  assign _0069_ = ~ div_valid;
  assign _0156_ = _0027_ & _0042_;
  assign _0159_ = _0566_ & _0044_;
  assign _0231_ = mult_en_internal_t0 & _0033_;
  assign _0234_ = { 1'h0, op_quotient_q_t0 } & _0067_;
  assign _0237_ = mult_valid_t0 & _0069_;
  assign _0157_ = _0558_ & _0041_;
  assign _0160_ = _0564_ & _0043_;
  assign _0232_ = div_en_internal_t0 & _0034_;
  assign _0235_ = { 1'h0, one_shift_t0 } & _0066_;
  assign _0238_ = div_valid_t0 & _0068_;
  assign _0158_ = _0027_ & _0558_;
  assign _0161_ = _0566_ & _0564_;
  assign _0233_ = mult_en_internal_t0 & div_en_internal_t0;
  assign _0236_ = { 1'h0, op_quotient_q_t0 } & { 1'h0, one_shift_t0 };
  assign _0239_ = mult_valid_t0 & div_valid_t0;
  assign _0348_ = _0156_ | _0157_;
  assign _0349_ = _0159_ | _0160_;
  assign _0404_ = _0231_ | _0232_;
  assign _0405_ = _0234_ | _0235_;
  assign _0406_ = _0237_ | _0238_;
  assign _0308_ = _0348_ | _0158_;
  assign _0310_ = _0349_ | _0161_;
  assign multdiv_en_t0 = _0404_ | _0233_;
  assign _0556_ = _0405_ | _0236_;
  assign valid_o_t0 = _0406_ | _0239_;
  assign _0307_ = _0026_ | _0557_;
  assign _0309_ = _0565_ | _0563_;
  assign _0092_ = | { _0567_, _0559_, _0557_ };
  assign \gen_mult_single_cycle.mult_state_d  = \gen_mult_single_cycle.mult_state_q  ? 1'h0 : _0000_;
  assign mult_hold = \gen_mult_single_cycle.mult_state_q  ? _0485_ : _0006_;
  assign mac_res_d = \gen_mult_single_cycle.mult_state_q  ? mac_res_ext[33:0] : _0002_;
  assign mult_valid = \gen_mult_single_cycle.mult_state_q  ? 1'h1 : _0008_;
  assign \gen_mult_single_cycle.summand2  = \gen_mult_single_cycle.mult_state_q  ? { accum[33], accum[33], accum[33], accum[33], accum[33], accum[33], accum[33], accum[33], accum[33], accum[33], accum[33], accum[33], accum[33], accum[33], accum[33], accum[33], imd_val_q_i[67:50] } : \gen_mult_single_cycle.mult2_res ;
  assign \gen_mult_single_cycle.summand1  = \gen_mult_single_cycle.mult_state_q  ? 34'h000000000 : { 18'h00000, \gen_mult_single_cycle.mult1_res [31:16] };
  assign \gen_mult_single_cycle.mult3_sign_b  = \gen_mult_single_cycle.mult_state_q  ? div_sign_b : 1'h0;
  assign \gen_mult_single_cycle.mult3_op_b  = \gen_mult_single_cycle.mult_state_q  ? op_b_i[31:16] : op_b_i[15:0];
  assign _0515_ = _0557_ ? { _0554_, 1'h1 } : { _0553_, 1'h1 };
  assign _0517_ = _0565_ ? { _0552_, 1'h1 } : { _0551_, 1'h1 };
  assign alu_operand_b_o = _0307_ ? _0515_ : _0517_;
  assign _0519_ = _0559_ ? 3'h5 : _0577_;
  assign _0521_ = _0557_ ? 3'h6 : _0519_;
  assign _0523_ = _0563_ ? 3'h3 : 3'h2;
  assign _0525_ = _0561_ ? _0004_ : 3'h0;
  assign _0527_ = _0309_ ? _0523_ : _0525_;
  assign md_state_d = _0092_ ? _0521_ : _0527_;
  assign _0529_ = _0559_ ? _0012_ : { 1'h0, next_remainder, _0570_ };
  assign _0531_ = _0557_ ? _0014_ : _0529_;
  assign _0533_ = _0561_ ? _0010_ : imd_val_q_i[67:34];
  assign _0535_ = _0563_ ? { 33'h000000000, op_numerator_q[31] } : _0533_;
  assign op_remainder_d = _0092_ ? _0531_ : _0535_;
  assign op_quotient_d = _0567_ ? next_quotient[31:0] : 32'd0;
  assign _0095_ = | { _0019_, div_en_internal_t0 };
  assign _0096_ = | { _0566_, div_en_internal_t0 };
  assign _0097_ = | { _0562_, _0541_, div_en_internal_t0 };
  assign _0345_ = { _0018_, div_en_internal } | { _0019_, div_en_internal_t0 };
  assign _0346_ = { _0565_, div_en_internal } | { _0566_, div_en_internal_t0 };
  assign _0347_ = { _0561_, _0540_, div_en_internal } | { _0562_, _0541_, div_en_internal_t0 };
  assign _0089_ = & _0345_;
  assign _0090_ = & _0346_;
  assign _0091_ = & _0347_;
  assign _0021_ = _0095_ & _0089_;
  assign _0023_ = _0096_ & _0090_;
  assign _0025_ = _0097_ & _0091_;
  assign _0105_ = | _0430_;
  wire [31:0] _1253_ = op_numerator_q_t0;
  assign _0537_ = _1253_[_0572_ +: 1];
  assign _0571_ = _0105_ | _0537_;
  assign _0101_ = | div_counter_q_t0;
  assign _0538_ = 32'd0 << div_counter_q;
  assign one_shift_t0 = { _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_ } | _0538_;
  assign _0429_ = div_counter_q | div_counter_q_t0;
  assign _0513_ = _0429_ - 5'h01;
  assign _0514_ = _0223_ - 5'h01;
  assign _0493_ = _0513_ ^ _0514_;
  assign _0430_ = _0493_ | div_counter_q_t0;
  assign _0584_ = imd_val_q_i_t0[65] | imd_val_q_i_t0[31];
  assign _0586_ = div_sign_a_t0 | div_sign_b_t0;
  assign _0539_ = ~ alu_adder_ext_i[32];
  assign _0542_ = div_counter_q == 5'h01;
  assign _0540_ = operator_i == 2'h2;
  assign _0544_ = _0546_ && equal_to_zero_i;
  assign _0546_ = ! data_ind_timing_i;
  assign \gen_mult_single_cycle.mult1_res  = $signed({ 18'h00000, op_a_i[15:0] }) * $signed({ 18'h00000, op_b_i[15:0] });
  assign \gen_mult_single_cycle.mult2_res  = $signed({ 18'h00000, op_a_i[15:0] }) * $signed({ div_sign_b, div_sign_b, div_sign_b, div_sign_b, div_sign_b, div_sign_b, div_sign_b, div_sign_b, div_sign_b, div_sign_b, div_sign_b, div_sign_b, div_sign_b, div_sign_b, div_sign_b, div_sign_b, div_sign_b, div_sign_b, op_b_i[31:16] });
  assign \gen_mult_single_cycle.mult3_res  = $signed({ div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, div_sign_a, op_a_i[31:16] }) * $signed({ \gen_mult_single_cycle.mult3_sign_b , \gen_mult_single_cycle.mult3_sign_b , \gen_mult_single_cycle.mult3_sign_b , \gen_mult_single_cycle.mult3_sign_b , \gen_mult_single_cycle.mult3_sign_b , \gen_mult_single_cycle.mult3_sign_b , \gen_mult_single_cycle.mult3_sign_b , \gen_mult_single_cycle.mult3_sign_b , \gen_mult_single_cycle.mult3_sign_b , \gen_mult_single_cycle.mult3_sign_b , \gen_mult_single_cycle.mult3_sign_b , \gen_mult_single_cycle.mult3_sign_b , \gen_mult_single_cycle.mult3_sign_b , \gen_mult_single_cycle.mult3_sign_b , \gen_mult_single_cycle.mult3_sign_b , \gen_mult_single_cycle.mult3_sign_b , \gen_mult_single_cycle.mult3_sign_b , \gen_mult_single_cycle.mult3_sign_b , \gen_mult_single_cycle.mult3_op_b  });
  assign signed_mult = | signed_mode_i;
  assign _0547_ = | operator_i;
  assign _0548_ = ~ mult_hold;
  assign _0549_ = ~ div_hold;
  assign _0485_ = ~ multdiv_ready_id_i;
  assign _0550_ = ~ div_by_zero_q;
  assign _0552_ = ~ op_a_i;
  assign _0551_ = ~ op_b_i;
  assign _0553_ = ~ imd_val_q_i[31:0];
  assign _0554_ = ~ imd_val_q_i[65:34];
  assign multdiv_en = mult_en_internal | div_en_internal;
  assign _0555_ = { 1'h0, op_quotient_q } | { 1'h0, one_shift };
  assign valid_o = mult_valid | div_valid;
  assign _0000_ = _0547_ ? 1'h1 : 1'h0;
  assign _0008_ = _0547_ ? 1'h0 : mult_en_i;
  assign _0002_ = _0547_ ? mac_res_ext[33:0] : { 2'h0, mac_res_ext[15:0], \gen_mult_single_cycle.mult1_res [15:0] };
  assign _0006_ = _0547_ ? 1'h0 : _0485_;
  assign _0014_ = _0540_ ? _0579_ : _0581_;
  assign _0012_ = _0540_ ? { 1'h0, next_quotient } : { 2'h0, next_remainder };
  assign _0010_ = _0540_ ? 34'h3ffffffff : { 2'h0, op_a_i };
  assign div_counter_d = _0028_ ? 5'h1f : _0572_;
  assign alu_operand_a_o = _0026_ ? { imd_val_q_i[65:34], 1'h1 } : 33'h000000001;
  assign _0557_ = md_state_q == 3'h5;
  assign _0559_ = md_state_q == 3'h4;
  assign _0561_ = ! md_state_q;
  assign div_hold = _0569_ ? _0485_ : 1'h0;
  assign div_valid = _0569_ ? 1'h1 : 1'h0;
  assign _0569_ = md_state_q == 3'h6;
  assign _0567_ = md_state_q == 3'h3;
  assign _0565_ = md_state_q == 3'h1;
  assign op_denominator_d = _0563_ ? _0575_ : imd_val_q_i[31:0];
  assign _0563_ = md_state_q == 3'h2;
  assign is_greater_equal = _0583_ ? imd_val_q_i[65] : _0539_;
  wire [31:0] _1254_ = op_numerator_q;
  assign _0570_ = _1254_[_0572_ +: 1];
  assign one_shift = 32'd1 << div_counter_q;
  assign _0572_ = div_counter_q - 5'h01;
  assign imd_val_d_o[67:34] = div_sel_i ? op_remainder_d : mac_res_d;
  assign multdiv_result_o = div_sel_i ? imd_val_q_i[65:34] : mac_res_d[31:0];
  assign next_remainder = is_greater_equal ? alu_adder_ext_i[32:1] : imd_val_q_i[65:34];
  assign next_quotient = is_greater_equal ? _0555_ : { 1'h0, op_quotient_q };
  assign _0004_ = _0544_ ? 3'h6 : 3'h1;
  assign _0573_ = div_sign_a ? alu_adder_i : op_a_i;
  assign _0575_ = div_sign_b ? alu_adder_i : op_b_i;
  assign _0577_ = _0542_ ? 3'h4 : 3'h3;
  assign _0579_ = div_change_sign ? { 2'h0, alu_adder_i } : imd_val_q_i[67:34];
  assign _0581_ = div_sign_a ? { 2'h0, alu_adder_i } : imd_val_q_i[67:34];
  assign _0583_ = imd_val_q_i[65] ^ imd_val_q_i[31];
  assign _0585_ = div_sign_a ^ div_sign_b;
  assign accum[32:0] = { accum[33], accum[33], accum[33], accum[33], accum[33], accum[33], accum[33], accum[33], accum[33], accum[33], accum[33], accum[33], accum[33], accum[33], accum[33], imd_val_q_i[67:50] };
  assign accum_t0[32:0] = { accum_t0[33], accum_t0[33], accum_t0[33], accum_t0[33], accum_t0[33], accum_t0[33], accum_t0[33], accum_t0[33], accum_t0[33], accum_t0[33], accum_t0[33], accum_t0[33], accum_t0[33], accum_t0[33], accum_t0[33], imd_val_q_i_t0[67:50] };
  assign imd_val_d_o[33:0] = { 2'h0, op_denominator_d };
  assign imd_val_d_o_t0[33:0] = { 2'h0, op_denominator_d_t0 };
  assign imd_val_we_o = { div_en_internal, multdiv_en };
  assign imd_val_we_o_t0 = { div_en_internal_t0, multdiv_en_t0 };
endmodule

module paramodauxy_ibex_prefetch_bufferBranchPredictor10 (clk_i, rst_ni, req_i, branch_i, branch_spec_i, predicted_branch_i, branch_mispredict_i, addr_i, ready_i, valid_o, rdata_o, addr_o, err_o, err_plus2_o, instr_req_o, instr_gnt_i, instr_addr_o, instr_rdata_i, instr_err_i, instr_pmp_err_i, instr_rvalid_i
, busy_o, valid_o_t0, req_i_t0, ready_i_t0, predicted_branch_i_t0, instr_rvalid_i_t0, instr_req_o_t0, instr_rdata_i_t0, instr_pmp_err_i_t0, instr_gnt_i_t0, instr_err_i_t0, instr_addr_o_t0, err_plus2_o_t0, err_o_t0, branch_spec_i_t0, branch_mispredict_i_t0, branch_i_t0, addr_o_t0, addr_i_t0, busy_o_t0, rdata_o_t0
);
  wire _000_;
  wire _001_;
  wire _002_;
  wire _003_;
  wire _004_;
  wire _005_;
  wire _006_;
  wire _007_;
  wire _008_;
  wire _009_;
  wire _010_;
  wire _011_;
  wire _012_;
  wire _013_;
  wire _014_;
  wire _015_;
  wire _016_;
  wire _017_;
  wire _018_;
  wire _019_;
  wire _020_;
  wire _021_;
  wire _022_;
  wire _023_;
  wire _024_;
  wire _025_;
  wire _026_;
  wire _027_;
  wire _028_;
  wire _029_;
  wire [31:0] _030_;
  wire [31:0] _031_;
  wire _032_;
  wire _033_;
  wire _034_;
  wire _035_;
  wire _036_;
  wire _037_;
  wire _038_;
  wire _039_;
  wire _040_;
  wire [1:0] _041_;
  wire [1:0] _042_;
  wire _043_;
  wire _044_;
  wire _045_;
  wire _046_;
  wire _047_;
  wire _048_;
  wire _049_;
  wire _050_;
  wire _051_;
  wire _052_;
  wire _053_;
  wire _054_;
  wire _055_;
  wire _056_;
  wire _057_;
  wire _058_;
  wire _059_;
  wire _060_;
  wire _061_;
  wire _062_;
  wire _063_;
  wire _064_;
  wire _065_;
  wire _066_;
  wire [1:0] _067_;
  wire [31:0] _068_;
  wire [31:0] _069_;
  wire [31:0] _070_;
  wire [31:0] _071_;
  wire [1:0] _072_;
  wire _073_;
  wire _074_;
  wire _075_;
  wire _076_;
  wire _077_;
  wire _078_;
  wire [31:0] _079_;
  wire [31:0] _080_;
  wire _081_;
  wire _082_;
  wire _083_;
  wire _084_;
  wire _085_;
  wire _086_;
  wire _087_;
  wire _088_;
  wire _089_;
  wire _090_;
  wire _091_;
  wire _092_;
  wire _093_;
  wire _094_;
  wire _095_;
  wire _096_;
  wire _097_;
  wire _098_;
  wire _099_;
  wire _100_;
  wire _101_;
  wire _102_;
  wire _103_;
  wire _104_;
  wire _105_;
  wire _106_;
  wire _107_;
  wire _108_;
  wire _109_;
  wire _110_;
  wire _111_;
  wire _112_;
  wire _113_;
  wire _114_;
  wire _115_;
  wire _116_;
  wire _117_;
  wire _118_;
  wire _119_;
  wire _120_;
  wire _121_;
  wire _122_;
  wire _123_;
  wire _124_;
  wire _125_;
  wire _126_;
  wire _127_;
  wire _128_;
  wire _129_;
  wire _130_;
  wire _131_;
  wire _132_;
  wire _133_;
  wire _134_;
  wire _135_;
  wire _136_;
  wire _137_;
  wire _138_;
  wire _139_;
  wire _140_;
  wire _141_;
  wire _142_;
  wire _143_;
  wire _144_;
  wire [31:0] _145_;
  wire [31:0] _146_;
  wire [31:0] _147_;
  wire [1:0] _148_;
  wire [1:0] _149_;
  wire [1:0] _150_;
  wire [29:0] _151_;
  wire [29:0] _152_;
  wire [29:0] _153_;
  wire _154_;
  wire _155_;
  wire _156_;
  wire _157_;
  wire _158_;
  wire _159_;
  wire _160_;
  wire _161_;
  wire _162_;
  wire [1:0] _163_;
  wire [1:0] _164_;
  wire [1:0] _165_;
  wire _166_;
  wire _167_;
  wire _168_;
  wire _169_;
  wire _170_;
  wire _171_;
  wire _172_;
  wire _173_;
  wire _174_;
  wire _175_;
  wire _176_;
  wire _177_;
  wire _178_;
  wire _179_;
  wire _180_;
  wire _181_;
  wire _182_;
  wire _183_;
  wire _184_;
  wire _185_;
  wire _186_;
  wire _187_;
  wire _188_;
  wire _189_;
  wire _190_;
  wire _191_;
  wire _192_;
  wire _193_;
  wire _194_;
  wire _195_;
  wire _196_;
  wire _197_;
  wire _198_;
  wire _199_;
  wire _200_;
  wire _201_;
  wire _202_;
  wire _203_;
  wire _204_;
  wire [1:0] _205_;
  wire [31:0] _206_;
  wire [31:0] _207_;
  wire [31:0] _208_;
  wire [31:0] _209_;
  wire [31:0] _210_;
  wire [31:0] _211_;
  wire [31:0] _212_;
  wire [31:0] _213_;
  wire [31:0] _214_;
  wire [31:0] _215_;
  wire [31:0] _216_;
  wire [31:0] _217_;
  wire [31:0] _218_;
  wire [31:0] _219_;
  wire [1:0] _220_;
  wire [1:0] _221_;
  wire [1:0] _222_;
  wire [1:0] _223_;
  wire [1:0] _224_;
  wire [1:0] _225_;
  wire [1:0] _226_;
  wire [1:0] _227_;
  wire [1:0] _228_;
  wire [31:0] _229_;
  wire [31:0] _230_;
  wire [31:0] _231_;
  wire [31:0] _232_;
  wire [31:0] _233_;
  wire _234_;
  wire _235_;
  wire _236_;
  wire _237_;
  wire _238_;
  wire _239_;
  wire _240_;
  wire _241_;
  wire _242_;
  wire _243_;
  wire _244_;
  wire _245_;
  wire _246_;
  wire _247_;
  wire _248_;
  wire _249_;
  wire _250_;
  wire _251_;
  wire _252_;
  wire _253_;
  wire _254_;
  wire _255_;
  wire [31:0] _256_;
  wire [31:0] _257_;
  wire [31:0] _258_;
  wire [31:0] _259_;
  wire [1:0] _260_;
  wire [1:0] _261_;
  wire [1:0] _262_;
  wire [1:0] _263_;
  wire [29:0] _264_;
  wire [29:0] _265_;
  wire [29:0] _266_;
  wire [29:0] _267_;
  wire [1:0] _268_;
  wire _269_;
  wire _270_;
  wire _271_;
  wire [1:0] _272_;
  wire _273_;
  wire _274_;
  wire _275_;
  wire _276_;
  wire _277_;
  wire _278_;
  wire _279_;
  wire _280_;
  wire _281_;
  wire _282_;
  wire _283_;
  wire _284_;
  wire _285_;
  wire _286_;
  wire [1:0] _287_;
  wire [31:0] _288_;
  wire [31:0] _289_;
  wire [31:0] _290_;
  wire [31:0] _291_;
  wire [31:0] _292_;
  wire [31:0] _293_;
  wire [31:0] _294_;
  wire [31:0] _295_;
  wire [31:0] _296_;
  wire [31:0] _297_;
  wire [31:0] _298_;
  wire [31:0] _299_;
  wire [31:0] _300_;
  wire [1:0] _301_;
  wire [1:0] _302_;
  wire [1:0] _303_;
  wire [1:0] _304_;
  wire [1:0] _305_;
  wire [31:0] _306_;
  wire [31:0] _307_;
  wire [31:0] _308_;
  wire [1:0] _309_;
  wire [29:0] _310_;
  wire [31:0] _311_;
  wire [31:0] _312_;
  wire [31:0] _313_;
  wire [1:0] _314_;
  wire [1:0] _315_;
  wire [1:0] _316_;
  wire [31:0] _317_;
  wire [31:0] _318_;
  wire _319_;
  wire _320_;
  wire [1:0] _321_;
  wire [1:0] _322_;
  wire _323_;
  wire _324_;
  wire _325_;
  wire _326_;
  wire _327_;
  wire _328_;
  wire _329_;
  wire _330_;
  wire _331_;
  wire _332_;
  wire _333_;
  wire _334_;
  wire [31:0] _335_;
  wire [31:0] _336_;
  wire [31:0] _337_;
  wire [31:0] _338_;
  wire [31:0] _339_;
  wire [31:0] _340_;
  wire [31:0] _341_;
  wire [31:0] _342_;
  input [31:0] addr_i;
  wire [31:0] addr_i;
  input [31:0] addr_i_t0;
  wire [31:0] addr_i_t0;
  wire [31:0] addr_next;
  wire [31:0] addr_next_t0;
  output [31:0] addr_o;
  wire [31:0] addr_o;
  output [31:0] addr_o_t0;
  wire [31:0] addr_o_t0;
  wire [1:0] branch_discard_n;
  wire [1:0] branch_discard_n_t0;
  reg [1:0] branch_discard_q;
  reg [1:0] branch_discard_q_t0;
  wire [1:0] branch_discard_s;
  wire [1:0] branch_discard_s_t0;
  input branch_i;
  wire branch_i;
  input branch_i_t0;
  wire branch_i_t0;
  input branch_mispredict_i;
  wire branch_mispredict_i;
  input branch_mispredict_i_t0;
  wire branch_mispredict_i_t0;
  wire branch_or_mispredict;
  wire branch_or_mispredict_t0;
  input branch_spec_i;
  wire branch_spec_i;
  input branch_spec_i_t0;
  wire branch_spec_i_t0;
  wire branch_suppress;
  wire branch_suppress_t0;
  output busy_o;
  wire busy_o;
  output busy_o_t0;
  wire busy_o_t0;
  input clk_i;
  wire clk_i;
  wire discard_req_d;
  wire discard_req_d_t0;
  reg discard_req_q;
  reg discard_req_q_t0;
  output err_o;
  wire err_o;
  output err_o_t0;
  wire err_o_t0;
  output err_plus2_o;
  wire err_plus2_o;
  output err_plus2_o_t0;
  wire err_plus2_o_t0;
  wire [31:0] fetch_addr_d;
  wire [31:0] fetch_addr_d_t0;
  wire fetch_addr_en;
  wire fetch_addr_en_t0;
  reg [31:0] fetch_addr_q;
  reg [31:0] fetch_addr_q_t0;
  wire [31:0] fifo_addr;
  wire [31:0] fifo_addr_t0;
  wire [1:0] fifo_busy;
  wire [1:0] fifo_busy_t0;
  wire fifo_ready;
  wire fifo_ready_t0;
  wire fifo_valid;
  wire fifo_valid_t0;
  wire gnt_or_pmp_err;
  wire gnt_or_pmp_err_t0;
  wire [31:0] instr_addr;
  output [31:0] instr_addr_o;
  wire [31:0] instr_addr_o;
  output [31:0] instr_addr_o_t0;
  wire [31:0] instr_addr_o_t0;
  wire [31:0] instr_addr_t0;
  input instr_err_i;
  wire instr_err_i;
  input instr_err_i_t0;
  wire instr_err_i_t0;
  input instr_gnt_i;
  wire instr_gnt_i;
  input instr_gnt_i_t0;
  wire instr_gnt_i_t0;
  wire instr_or_pmp_err;
  wire instr_or_pmp_err_t0;
  input instr_pmp_err_i;
  wire instr_pmp_err_i;
  input instr_pmp_err_i_t0;
  wire instr_pmp_err_i_t0;
  input [31:0] instr_rdata_i;
  wire [31:0] instr_rdata_i;
  input [31:0] instr_rdata_i_t0;
  wire [31:0] instr_rdata_i_t0;
  output instr_req_o;
  wire instr_req_o;
  output instr_req_o_t0;
  wire instr_req_o_t0;
  input instr_rvalid_i;
  wire instr_rvalid_i;
  input instr_rvalid_i_t0;
  wire instr_rvalid_i_t0;
  input predicted_branch_i;
  wire predicted_branch_i;
  input predicted_branch_i_t0;
  wire predicted_branch_i_t0;
  output [31:0] rdata_o;
  wire [31:0] rdata_o;
  output [31:0] rdata_o_t0;
  wire [31:0] rdata_o_t0;
  wire [1:0] rdata_outstanding_n;
  wire [1:0] rdata_outstanding_n_t0;
  reg [1:0] rdata_outstanding_q;
  reg [1:0] rdata_outstanding_q_t0;
  wire [1:0] rdata_outstanding_s;
  wire [1:0] rdata_outstanding_s_t0;
  wire [1:0] rdata_pmp_err_n;
  wire [1:0] rdata_pmp_err_n_t0;
  reg [1:0] rdata_pmp_err_q;
  reg [1:0] rdata_pmp_err_q_t0;
  wire [1:0] rdata_pmp_err_s;
  wire [1:0] rdata_pmp_err_s_t0;
  input ready_i;
  wire ready_i;
  input ready_i_t0;
  wire ready_i_t0;
  input req_i;
  wire req_i;
  input req_i_t0;
  wire req_i_t0;
  input rst_ni;
  wire rst_ni;
  wire rvalid_or_pmp_err;
  wire rvalid_or_pmp_err_t0;
  wire stored_addr_en;
  wire stored_addr_en_t0;
  reg [31:0] stored_addr_q;
  reg [31:0] stored_addr_q_t0;
  wire valid_new_req;
  wire valid_new_req_t0;
  output valid_o;
  wire valid_o;
  output valid_o_t0;
  wire valid_o_t0;
  wire valid_raw;
  wire valid_raw_t0;
  wire valid_req_d;
  wire valid_req_d_t0;
  reg valid_req_q;
  reg valid_req_q_t0;
  assign fetch_addr_d = _337_ + { 29'h00000000, _004_, 2'h0 };
  assign branch_suppress = branch_spec_i & _037_;
  assign _000_ = _319_ & req_i;
  assign _002_ = _000_ & _323_;
  assign valid_new_req = _002_ & _060_;
  assign rvalid_or_pmp_err = rdata_outstanding_q[0] & _325_;
  assign valid_req_d = instr_req_o & _320_;
  assign discard_req_d = valid_req_q & _327_;
  assign stored_addr_en = _004_ & _320_;
  assign _004_ = valid_new_req & _045_;
  assign _010_ = branch_or_mispredict & rdata_outstanding_q[0];
  assign _012_ = instr_req_o & _053_;
  assign _014_ = _012_ & instr_pmp_err_i;
  assign _016_ = _006_ & rdata_outstanding_q[0];
  assign _006_ = instr_req_o & gnt_or_pmp_err;
  assign _008_ = _006_ & discard_req_d;
  assign _018_ = _008_ & rdata_outstanding_q[0];
  assign _020_ = branch_or_mispredict & rdata_outstanding_q[1];
  assign _022_ = instr_req_o & _060_;
  assign _024_ = _022_ & instr_pmp_err_i;
  assign _026_ = _024_ & rdata_outstanding_q[0];
  assign fifo_valid = rvalid_or_pmp_err & _057_;
  assign valid_o = valid_raw & _038_;
  assign _030_ = ~ _338_;
  assign _031_ = ~ { 29'h00000000, _005_, 2'h0 };
  assign _079_ = _337_ & _030_;
  assign _080_ = { 29'h00000000, _004_, 2'h0 } & _031_;
  assign _317_ = _079_ + _080_;
  assign _231_ = _337_ | _338_;
  assign _232_ = { 29'h00000000, _004_, 2'h0 } | { 29'h00000000, _005_, 2'h0 };
  assign _318_ = _231_ + _232_;
  assign _307_ = _317_ ^ _318_;
  assign _233_ = _307_ | _338_;
  assign fetch_addr_d_t0 = _233_ | { 29'h00000000, _005_, 2'h0 };
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) valid_req_q_t0 <= 1'h0;
    else valid_req_q_t0 <= valid_req_d_t0;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) discard_req_q_t0 <= 1'h0;
    else discard_req_q_t0 <= discard_req_d_t0;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) rdata_outstanding_q_t0 <= 2'h0;
    else rdata_outstanding_q_t0 <= rdata_outstanding_s_t0;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) branch_discard_q_t0 <= 2'h0;
    else branch_discard_q_t0 <= branch_discard_s_t0;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) rdata_pmp_err_q_t0 <= 2'h0;
    else rdata_pmp_err_q_t0 <= rdata_pmp_err_s_t0;
  assign _081_ = branch_spec_i_t0 & _037_;
  assign _084_ = branch_suppress_t0 & req_i;
  assign _087_ = _001_ & _323_;
  assign _090_ = _003_ & _060_;
  assign _093_ = rdata_outstanding_q_t0[0] & _325_;
  assign _096_ = instr_req_o_t0 & _320_;
  assign _099_ = valid_req_q_t0 & _327_;
  assign _102_ = _005_ & _320_;
  assign _108_ = branch_or_mispredict_t0 & rdata_outstanding_q[0];
  assign _111_ = instr_req_o_t0 & _053_;
  assign _114_ = _013_ & instr_pmp_err_i;
  assign _117_ = _007_ & rdata_outstanding_q[0];
  assign _120_ = instr_req_o_t0 & gnt_or_pmp_err;
  assign _121_ = _007_ & discard_req_d;
  assign _124_ = _009_ & rdata_outstanding_q[0];
  assign _127_ = branch_or_mispredict_t0 & rdata_outstanding_q[1];
  assign _130_ = instr_req_o_t0 & _060_;
  assign _133_ = _023_ & instr_pmp_err_i;
  assign _136_ = _025_ & rdata_outstanding_q[0];
  assign _139_ = rvalid_or_pmp_err_t0 & _057_;
  assign _142_ = valid_raw_t0 & _038_;
  assign _082_ = branch_i_t0 & branch_spec_i;
  assign _085_ = req_i_t0 & _319_;
  assign _088_ = _324_ & _000_;
  assign _091_ = rdata_outstanding_q_t0[1] & _002_;
  assign _094_ = _326_ & rdata_outstanding_q[0];
  assign _100_ = _328_ & valid_req_q;
  assign _103_ = gnt_or_pmp_err_t0 & _004_;
  assign _106_ = valid_req_q_t0 & valid_new_req;
  assign _109_ = rdata_outstanding_q_t0[0] & branch_or_mispredict;
  assign _112_ = rdata_outstanding_q_t0[0] & instr_req_o;
  assign _115_ = instr_pmp_err_i_t0 & _012_;
  assign _118_ = rdata_outstanding_q_t0[0] & _006_;
  assign _097_ = gnt_or_pmp_err_t0 & instr_req_o;
  assign _122_ = discard_req_d_t0 & _006_;
  assign _125_ = rdata_outstanding_q_t0[0] & _008_;
  assign _128_ = rdata_outstanding_q_t0[1] & branch_or_mispredict;
  assign _131_ = rdata_outstanding_q_t0[1] & instr_req_o;
  assign _134_ = instr_pmp_err_i_t0 & _022_;
  assign _137_ = rdata_outstanding_q_t0[0] & _024_;
  assign _140_ = branch_discard_q_t0[0] & rvalid_or_pmp_err;
  assign _143_ = branch_mispredict_i_t0 & valid_raw;
  assign _083_ = branch_spec_i_t0 & branch_i_t0;
  assign _086_ = branch_suppress_t0 & req_i_t0;
  assign _089_ = _001_ & _324_;
  assign _092_ = _003_ & rdata_outstanding_q_t0[1];
  assign _095_ = rdata_outstanding_q_t0[0] & _326_;
  assign _101_ = valid_req_q_t0 & _328_;
  assign _104_ = _005_ & gnt_or_pmp_err_t0;
  assign _110_ = branch_or_mispredict_t0 & rdata_outstanding_q_t0[0];
  assign _113_ = instr_req_o_t0 & rdata_outstanding_q_t0[0];
  assign _116_ = _013_ & instr_pmp_err_i_t0;
  assign _098_ = instr_req_o_t0 & gnt_or_pmp_err_t0;
  assign _123_ = _007_ & discard_req_d_t0;
  assign _126_ = _009_ & rdata_outstanding_q_t0[0];
  assign _129_ = branch_or_mispredict_t0 & rdata_outstanding_q_t0[1];
  assign _132_ = instr_req_o_t0 & rdata_outstanding_q_t0[1];
  assign _135_ = _023_ & instr_pmp_err_i_t0;
  assign _138_ = _025_ & rdata_outstanding_q_t0[0];
  assign _141_ = rvalid_or_pmp_err_t0 & branch_discard_q_t0[0];
  assign _144_ = valid_raw_t0 & branch_mispredict_i_t0;
  assign _234_ = _081_ | _082_;
  assign _235_ = _084_ | _085_;
  assign _236_ = _087_ | _088_;
  assign _237_ = _090_ | _091_;
  assign _238_ = _093_ | _094_;
  assign _239_ = _096_ | _097_;
  assign _240_ = _099_ | _100_;
  assign _241_ = _102_ | _103_;
  assign _242_ = _105_ | _106_;
  assign _243_ = _108_ | _109_;
  assign _244_ = _111_ | _112_;
  assign _245_ = _114_ | _115_;
  assign _246_ = _117_ | _118_;
  assign _247_ = _120_ | _097_;
  assign _248_ = _121_ | _122_;
  assign _249_ = _124_ | _125_;
  assign _250_ = _127_ | _128_;
  assign _251_ = _130_ | _131_;
  assign _252_ = _133_ | _134_;
  assign _253_ = _136_ | _137_;
  assign _254_ = _139_ | _140_;
  assign _255_ = _142_ | _143_;
  assign branch_suppress_t0 = _234_ | _083_;
  assign _001_ = _235_ | _086_;
  assign _003_ = _236_ | _089_;
  assign valid_new_req_t0 = _237_ | _092_;
  assign rvalid_or_pmp_err_t0 = _238_ | _095_;
  assign valid_req_d_t0 = _239_ | _098_;
  assign discard_req_d_t0 = _240_ | _101_;
  assign stored_addr_en_t0 = _241_ | _104_;
  assign _005_ = _242_ | _107_;
  assign _011_ = _243_ | _110_;
  assign _013_ = _244_ | _113_;
  assign _015_ = _245_ | _116_;
  assign _017_ = _246_ | _119_;
  assign _007_ = _247_ | _098_;
  assign _009_ = _248_ | _123_;
  assign _019_ = _249_ | _126_;
  assign _021_ = _250_ | _129_;
  assign _023_ = _251_ | _132_;
  assign _025_ = _252_ | _135_;
  assign _027_ = _253_ | _138_;
  assign fifo_valid_t0 = _254_ | _141_;
  assign valid_o_t0 = _255_ | _144_;
  assign _308_ = fetch_addr_d ^ fetch_addr_q;
  assign _309_ = _341_[1:0] ^ stored_addr_q[1:0];
  assign _310_ = instr_addr[31:2] ^ stored_addr_q[31:2];
  assign _032_ = ~ fetch_addr_en;
  assign _033_ = ~ _028_;
  assign _034_ = ~ stored_addr_en;
  assign _256_ = fetch_addr_d_t0 | fetch_addr_q_t0;
  assign _260_ = _342_[1:0] | stored_addr_q_t0[1:0];
  assign _264_ = instr_addr_t0[31:2] | stored_addr_q_t0[31:2];
  assign _257_ = _308_ | _256_;
  assign _261_ = _309_ | _260_;
  assign _265_ = _310_ | _264_;
  assign _145_ = { fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en } & fetch_addr_d_t0;
  assign _148_ = { _028_, _028_ } & _342_[1:0];
  assign _151_ = { stored_addr_en, stored_addr_en, stored_addr_en, stored_addr_en, stored_addr_en, stored_addr_en, stored_addr_en, stored_addr_en, stored_addr_en, stored_addr_en, stored_addr_en, stored_addr_en, stored_addr_en, stored_addr_en, stored_addr_en, stored_addr_en, stored_addr_en, stored_addr_en, stored_addr_en, stored_addr_en, stored_addr_en, stored_addr_en, stored_addr_en, stored_addr_en, stored_addr_en, stored_addr_en, stored_addr_en, stored_addr_en, stored_addr_en, stored_addr_en } & instr_addr_t0[31:2];
  assign _146_ = { _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_ } & fetch_addr_q_t0;
  assign _149_ = { _033_, _033_ } & stored_addr_q_t0[1:0];
  assign _152_ = { _034_, _034_, _034_, _034_, _034_, _034_, _034_, _034_, _034_, _034_, _034_, _034_, _034_, _034_, _034_, _034_, _034_, _034_, _034_, _034_, _034_, _034_, _034_, _034_, _034_, _034_, _034_, _034_, _034_, _034_ } & stored_addr_q_t0[31:2];
  assign _147_ = _257_ & fetch_addr_en_t0;
  assign _150_ = _261_ & _029_;
  assign _153_ = _265_ & stored_addr_en_t0;
  assign _258_ = _145_ | _146_;
  assign _262_ = _148_ | _149_;
  assign _266_ = _151_ | _152_;
  assign _259_ = _258_ | _147_;
  assign _263_ = _262_ | _150_;
  assign _267_ = _266_ | _153_;
  always_ff @(posedge clk_i)
    fetch_addr_q_t0 <= _259_;
  always_ff @(posedge clk_i)
    stored_addr_q_t0[1:0] <= _263_;
  always_ff @(posedge clk_i)
    stored_addr_q_t0[31:2] <= _267_;
  always_ff @(posedge clk_i)
    if (fetch_addr_en) fetch_addr_q <= fetch_addr_d;
  always_ff @(posedge clk_i)
    if (_028_) stored_addr_q[1:0] <= _341_[1:0];
  always_ff @(posedge clk_i)
    if (stored_addr_en) stored_addr_q[31:2] <= instr_addr[31:2];
  assign _077_ = | rdata_outstanding_q_t0;
  assign _067_ = ~ rdata_outstanding_q_t0;
  assign _205_ = rdata_outstanding_q & _067_;
  assign _078_ = ! _205_;
  assign _334_ = _078_ & _077_;
  assign _068_ = ~ { branch_mispredict_i, branch_mispredict_i, branch_mispredict_i, branch_mispredict_i, branch_mispredict_i, branch_mispredict_i, branch_mispredict_i, branch_mispredict_i, branch_mispredict_i, branch_mispredict_i, branch_mispredict_i, branch_mispredict_i, branch_mispredict_i, branch_mispredict_i, branch_mispredict_i, branch_mispredict_i, branch_mispredict_i, branch_mispredict_i, branch_mispredict_i, branch_mispredict_i, branch_mispredict_i, branch_mispredict_i, branch_mispredict_i, branch_mispredict_i, branch_mispredict_i, branch_mispredict_i, branch_mispredict_i, branch_mispredict_i, branch_mispredict_i, branch_mispredict_i, branch_mispredict_i, branch_mispredict_i };
  assign _070_ = ~ { branch_spec_i, branch_spec_i, branch_spec_i, branch_spec_i, branch_spec_i, branch_spec_i, branch_spec_i, branch_spec_i, branch_spec_i, branch_spec_i, branch_spec_i, branch_spec_i, branch_spec_i, branch_spec_i, branch_spec_i, branch_spec_i, branch_spec_i, branch_spec_i, branch_spec_i, branch_spec_i, branch_spec_i, branch_spec_i, branch_spec_i, branch_spec_i, branch_spec_i, branch_spec_i, branch_spec_i, branch_spec_i, branch_spec_i, branch_spec_i, branch_spec_i, branch_spec_i };
  assign _071_ = ~ { valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q };
  assign _072_ = ~ { rvalid_or_pmp_err, rvalid_or_pmp_err };
  assign _069_ = ~ { branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i };
  assign _291_ = { branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0 } | _069_;
  assign _288_ = { branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0 } | _068_;
  assign _295_ = { branch_spec_i_t0, branch_spec_i_t0, branch_spec_i_t0, branch_spec_i_t0, branch_spec_i_t0, branch_spec_i_t0, branch_spec_i_t0, branch_spec_i_t0, branch_spec_i_t0, branch_spec_i_t0, branch_spec_i_t0, branch_spec_i_t0, branch_spec_i_t0, branch_spec_i_t0, branch_spec_i_t0, branch_spec_i_t0, branch_spec_i_t0, branch_spec_i_t0, branch_spec_i_t0, branch_spec_i_t0, branch_spec_i_t0, branch_spec_i_t0, branch_spec_i_t0, branch_spec_i_t0, branch_spec_i_t0, branch_spec_i_t0, branch_spec_i_t0, branch_spec_i_t0, branch_spec_i_t0, branch_spec_i_t0, branch_spec_i_t0, branch_spec_i_t0 } | _070_;
  assign _298_ = { valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0 } | _071_;
  assign _301_ = { rvalid_or_pmp_err_t0, rvalid_or_pmp_err_t0 } | _072_;
  assign _289_ = { branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0 } | { branch_mispredict_i, branch_mispredict_i, branch_mispredict_i, branch_mispredict_i, branch_mispredict_i, branch_mispredict_i, branch_mispredict_i, branch_mispredict_i, branch_mispredict_i, branch_mispredict_i, branch_mispredict_i, branch_mispredict_i, branch_mispredict_i, branch_mispredict_i, branch_mispredict_i, branch_mispredict_i, branch_mispredict_i, branch_mispredict_i, branch_mispredict_i, branch_mispredict_i, branch_mispredict_i, branch_mispredict_i, branch_mispredict_i, branch_mispredict_i, branch_mispredict_i, branch_mispredict_i, branch_mispredict_i, branch_mispredict_i, branch_mispredict_i, branch_mispredict_i, branch_mispredict_i, branch_mispredict_i };
  assign _296_ = { branch_spec_i_t0, branch_spec_i_t0, branch_spec_i_t0, branch_spec_i_t0, branch_spec_i_t0, branch_spec_i_t0, branch_spec_i_t0, branch_spec_i_t0, branch_spec_i_t0, branch_spec_i_t0, branch_spec_i_t0, branch_spec_i_t0, branch_spec_i_t0, branch_spec_i_t0, branch_spec_i_t0, branch_spec_i_t0, branch_spec_i_t0, branch_spec_i_t0, branch_spec_i_t0, branch_spec_i_t0, branch_spec_i_t0, branch_spec_i_t0, branch_spec_i_t0, branch_spec_i_t0, branch_spec_i_t0, branch_spec_i_t0, branch_spec_i_t0, branch_spec_i_t0, branch_spec_i_t0, branch_spec_i_t0, branch_spec_i_t0, branch_spec_i_t0 } | { branch_spec_i, branch_spec_i, branch_spec_i, branch_spec_i, branch_spec_i, branch_spec_i, branch_spec_i, branch_spec_i, branch_spec_i, branch_spec_i, branch_spec_i, branch_spec_i, branch_spec_i, branch_spec_i, branch_spec_i, branch_spec_i, branch_spec_i, branch_spec_i, branch_spec_i, branch_spec_i, branch_spec_i, branch_spec_i, branch_spec_i, branch_spec_i, branch_spec_i, branch_spec_i, branch_spec_i, branch_spec_i, branch_spec_i, branch_spec_i, branch_spec_i, branch_spec_i };
  assign _299_ = { valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0 } | { valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q };
  assign _302_ = { rvalid_or_pmp_err_t0, rvalid_or_pmp_err_t0 } | { rvalid_or_pmp_err, rvalid_or_pmp_err };
  assign _292_ = { branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0 } | { branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i };
  assign _206_ = { fetch_addr_q_t0[31:2], 2'h0 } & _288_;
  assign _209_ = _336_ & _291_;
  assign _212_ = fetch_addr_q_t0 & _288_;
  assign _214_ = _340_ & _295_;
  assign _217_ = _342_ & _298_;
  assign _220_ = rdata_outstanding_n_t0 & _301_;
  assign _223_ = branch_discard_n_t0 & _301_;
  assign _226_ = rdata_pmp_err_n_t0 & _301_;
  assign _229_ = 32'd0 & _291_;
  assign _207_ = 32'd0 & _289_;
  assign _215_ = addr_i_t0 & _296_;
  assign _218_ = stored_addr_q_t0 & _299_;
  assign _221_ = { 1'h0, rdata_outstanding_n_t0[1] } & _302_;
  assign _224_ = { 1'h0, branch_discard_n_t0[1] } & _302_;
  assign _227_ = { 1'h0, rdata_pmp_err_n_t0[1] } & _302_;
  assign _210_ = addr_i_t0 & _292_;
  assign _290_ = _206_ | _207_;
  assign _293_ = _209_ | _210_;
  assign _294_ = _212_ | _207_;
  assign _297_ = _214_ | _215_;
  assign _300_ = _217_ | _218_;
  assign _303_ = _220_ | _221_;
  assign _304_ = _223_ | _224_;
  assign _305_ = _226_ | _227_;
  assign _306_ = _229_ | _210_;
  assign _311_ = _335_ ^ addr_i;
  assign _312_ = _339_ ^ addr_i;
  assign _313_ = _341_ ^ stored_addr_q;
  assign _314_ = rdata_outstanding_n ^ { 1'h0, rdata_outstanding_n[1] };
  assign _315_ = branch_discard_n ^ { 1'h0, branch_discard_n[1] };
  assign _316_ = rdata_pmp_err_n ^ { 1'h0, rdata_pmp_err_n[1] };
  assign _208_ = { branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0 } & { fetch_addr_q[31:2], 2'h0 };
  assign _211_ = { branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0 } & _311_;
  assign _213_ = { branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0, branch_mispredict_i_t0 } & fetch_addr_q;
  assign _216_ = { branch_spec_i_t0, branch_spec_i_t0, branch_spec_i_t0, branch_spec_i_t0, branch_spec_i_t0, branch_spec_i_t0, branch_spec_i_t0, branch_spec_i_t0, branch_spec_i_t0, branch_spec_i_t0, branch_spec_i_t0, branch_spec_i_t0, branch_spec_i_t0, branch_spec_i_t0, branch_spec_i_t0, branch_spec_i_t0, branch_spec_i_t0, branch_spec_i_t0, branch_spec_i_t0, branch_spec_i_t0, branch_spec_i_t0, branch_spec_i_t0, branch_spec_i_t0, branch_spec_i_t0, branch_spec_i_t0, branch_spec_i_t0, branch_spec_i_t0, branch_spec_i_t0, branch_spec_i_t0, branch_spec_i_t0, branch_spec_i_t0, branch_spec_i_t0 } & _312_;
  assign _219_ = { valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0 } & _313_;
  assign _222_ = { rvalid_or_pmp_err_t0, rvalid_or_pmp_err_t0 } & _314_;
  assign _225_ = { rvalid_or_pmp_err_t0, rvalid_or_pmp_err_t0 } & _315_;
  assign _228_ = { rvalid_or_pmp_err_t0, rvalid_or_pmp_err_t0 } & _316_;
  assign _230_ = { branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0 } & addr_i;
  assign _336_ = _208_ | _290_;
  assign _338_ = _211_ | _293_;
  assign _340_ = _213_ | _294_;
  assign _342_ = _216_ | _297_;
  assign instr_addr_t0 = _219_ | _300_;
  assign rdata_outstanding_s_t0 = _222_ | _303_;
  assign branch_discard_s_t0 = _225_ | _304_;
  assign rdata_pmp_err_s_t0 = _228_ | _305_;
  assign fifo_addr_t0 = _230_ | _306_;
  assign _028_ = & { _045_, stored_addr_en };
  assign _035_ = ~ _333_;
  assign _037_ = ~ branch_i;
  assign _039_ = ~ instr_err_i;
  assign _041_ = ~ fifo_busy;
  assign _045_ = ~ valid_req_q;
  assign _047_ = ~ instr_gnt_i;
  assign _049_ = ~ instr_rvalid_i;
  assign _044_ = ~ branch_or_mispredict;
  assign _052_ = ~ _006_;
  assign _054_ = ~ _008_;
  assign _056_ = ~ _329_;
  assign _058_ = ~ _014_;
  assign _059_ = ~ _016_;
  assign _061_ = ~ _018_;
  assign _063_ = ~ _331_;
  assign _065_ = ~ _026_;
  assign _036_ = ~ instr_req_o;
  assign _038_ = ~ branch_mispredict_i;
  assign _042_ = ~ { rdata_outstanding_q[0], rdata_outstanding_q[1] };
  assign _046_ = ~ valid_new_req;
  assign _048_ = ~ instr_pmp_err_i;
  assign _050_ = ~ discard_req_q;
  assign _051_ = ~ _004_;
  assign _053_ = ~ rdata_outstanding_q[0];
  assign _055_ = ~ _010_;
  assign _057_ = ~ branch_discard_q[0];
  assign _040_ = ~ rdata_pmp_err_q[0];
  assign _060_ = ~ rdata_outstanding_q[1];
  assign _062_ = ~ _020_;
  assign _064_ = ~ branch_discard_q[1];
  assign _066_ = ~ rdata_pmp_err_q[1];
  assign _154_ = _334_ & _036_;
  assign _157_ = branch_i_t0 & _038_;
  assign _160_ = instr_err_i_t0 & _040_;
  assign _163_ = fifo_busy_t0 & _042_;
  assign _166_ = fifo_ready_t0 & _044_;
  assign _169_ = valid_req_q_t0 & _046_;
  assign _170_ = instr_gnt_i_t0 & _048_;
  assign _173_ = instr_rvalid_i_t0 & _040_;
  assign _176_ = branch_or_mispredict_t0 & _050_;
  assign _179_ = branch_or_mispredict_t0 & _051_;
  assign _182_ = _007_ & _053_;
  assign _184_ = _009_ & _055_;
  assign _187_ = _330_ & _057_;
  assign _190_ = _015_ & _040_;
  assign _193_ = _017_ & _060_;
  assign _196_ = _019_ & _062_;
  assign _199_ = _332_ & _064_;
  assign _202_ = _027_ & _066_;
  assign _155_ = instr_req_o_t0 & _035_;
  assign _158_ = branch_mispredict_i_t0 & _037_;
  assign _161_ = rdata_pmp_err_q_t0[0] & _039_;
  assign _164_ = { rdata_outstanding_q_t0[0], rdata_outstanding_q_t0[1] } & _041_;
  assign _167_ = branch_or_mispredict_t0 & _043_;
  assign _105_ = valid_new_req_t0 & _045_;
  assign _171_ = instr_pmp_err_i_t0 & _047_;
  assign _174_ = rdata_pmp_err_q_t0[0] & _049_;
  assign _177_ = discard_req_q_t0 & _044_;
  assign _180_ = _005_ & _044_;
  assign _183_ = rdata_outstanding_q_t0[0] & _052_;
  assign _185_ = _011_ & _054_;
  assign _188_ = branch_discard_q_t0[0] & _056_;
  assign _191_ = rdata_pmp_err_q_t0[0] & _058_;
  assign _194_ = rdata_outstanding_q_t0[1] & _059_;
  assign _197_ = _021_ & _061_;
  assign _200_ = branch_discard_q_t0[1] & _063_;
  assign _203_ = rdata_pmp_err_q_t0[1] & _065_;
  assign _156_ = _334_ & instr_req_o_t0;
  assign _159_ = branch_i_t0 & branch_mispredict_i_t0;
  assign _162_ = instr_err_i_t0 & rdata_pmp_err_q_t0[0];
  assign _165_ = fifo_busy_t0 & { rdata_outstanding_q_t0[0], rdata_outstanding_q_t0[1] };
  assign _168_ = fifo_ready_t0 & branch_or_mispredict_t0;
  assign _107_ = valid_req_q_t0 & valid_new_req_t0;
  assign _172_ = instr_gnt_i_t0 & instr_pmp_err_i_t0;
  assign _175_ = instr_rvalid_i_t0 & rdata_pmp_err_q_t0[0];
  assign _178_ = branch_or_mispredict_t0 & discard_req_q_t0;
  assign _181_ = branch_or_mispredict_t0 & _005_;
  assign _119_ = _007_ & rdata_outstanding_q_t0[0];
  assign _186_ = _009_ & _011_;
  assign _189_ = _330_ & branch_discard_q_t0[0];
  assign _192_ = _015_ & rdata_pmp_err_q_t0[0];
  assign _195_ = _017_ & rdata_outstanding_q_t0[1];
  assign _198_ = _019_ & _021_;
  assign _201_ = _332_ & branch_discard_q_t0[1];
  assign _204_ = _027_ & rdata_pmp_err_q_t0[1];
  assign _269_ = _154_ | _155_;
  assign _270_ = _157_ | _158_;
  assign _271_ = _160_ | _161_;
  assign _272_ = _163_ | _164_;
  assign _273_ = _166_ | _167_;
  assign _274_ = _169_ | _105_;
  assign _275_ = _170_ | _171_;
  assign _276_ = _173_ | _174_;
  assign _277_ = _176_ | _177_;
  assign _278_ = _179_ | _180_;
  assign _279_ = _182_ | _183_;
  assign _280_ = _184_ | _185_;
  assign _281_ = _187_ | _188_;
  assign _282_ = _190_ | _191_;
  assign _283_ = _193_ | _194_;
  assign _284_ = _196_ | _197_;
  assign _285_ = _199_ | _200_;
  assign _286_ = _202_ | _203_;
  assign busy_o_t0 = _269_ | _156_;
  assign branch_or_mispredict_t0 = _270_ | _159_;
  assign instr_or_pmp_err_t0 = _271_ | _162_;
  assign _322_ = _272_ | _165_;
  assign _324_ = _273_ | _168_;
  assign instr_req_o_t0 = _274_ | _107_;
  assign gnt_or_pmp_err_t0 = _275_ | _172_;
  assign _326_ = _276_ | _175_;
  assign _328_ = _277_ | _178_;
  assign fetch_addr_en_t0 = _278_ | _181_;
  assign rdata_outstanding_n_t0[0] = _279_ | _119_;
  assign _330_ = _280_ | _186_;
  assign branch_discard_n_t0[0] = _281_ | _189_;
  assign rdata_pmp_err_n_t0[0] = _282_ | _192_;
  assign rdata_outstanding_n_t0[1] = _283_ | _195_;
  assign _332_ = _284_ | _198_;
  assign branch_discard_n_t0[1] = _285_ | _201_;
  assign rdata_pmp_err_n_t0[1] = _286_ | _204_;
  assign _075_ = | { valid_req_q_t0, stored_addr_en_t0 };
  assign _076_ = | _322_;
  assign _268_ = { _045_, stored_addr_en } | { valid_req_q_t0, stored_addr_en_t0 };
  assign _287_ = _321_ | _322_;
  assign _073_ = & _268_;
  assign _074_ = & _287_;
  assign _029_ = _075_ & _073_;
  assign fifo_ready_t0 = _076_ & _074_;
  assign fifo_ready = ! _043_;
  assign _319_ = ~ branch_suppress;
  assign _320_ = ~ gnt_or_pmp_err;
  assign busy_o = _333_ | instr_req_o;
  assign branch_or_mispredict = branch_i | branch_mispredict_i;
  assign instr_or_pmp_err = instr_err_i | rdata_pmp_err_q[0];
  assign _321_ = fifo_busy | { rdata_outstanding_q[0], rdata_outstanding_q[1] };
  assign _323_ = fifo_ready | branch_or_mispredict;
  assign instr_req_o = valid_req_q | valid_new_req;
  assign gnt_or_pmp_err = instr_gnt_i | instr_pmp_err_i;
  assign _325_ = instr_rvalid_i | rdata_pmp_err_q[0];
  assign _327_ = branch_or_mispredict | discard_req_q;
  assign fetch_addr_en = branch_or_mispredict | _004_;
  assign rdata_outstanding_n[0] = _006_ | rdata_outstanding_q[0];
  assign _329_ = _008_ | _010_;
  assign branch_discard_n[0] = _329_ | branch_discard_q[0];
  assign rdata_pmp_err_n[0] = _014_ | rdata_pmp_err_q[0];
  assign rdata_outstanding_n[1] = _016_ | rdata_outstanding_q[1];
  assign _331_ = _018_ | _020_;
  assign branch_discard_n[1] = _331_ | branch_discard_q[1];
  assign rdata_pmp_err_n[1] = _026_ | rdata_pmp_err_q[1];
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) valid_req_q <= 1'h0;
    else valid_req_q <= valid_req_d;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) discard_req_q <= 1'h0;
    else discard_req_q <= discard_req_d;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) rdata_outstanding_q <= 2'h0;
    else rdata_outstanding_q <= rdata_outstanding_s;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) branch_discard_q <= 2'h0;
    else branch_discard_q <= branch_discard_s;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) rdata_pmp_err_q <= 2'h0;
    else rdata_pmp_err_q <= rdata_pmp_err_s;
  assign _043_ = & _321_;
  assign _333_ = | rdata_outstanding_q;
  assign _335_ = branch_mispredict_i ? 32'd0 : { fetch_addr_q[31:2], 2'h0 };
  assign _337_ = branch_i ? addr_i : _335_;
  assign _339_ = branch_mispredict_i ? 32'd0 : fetch_addr_q;
  assign _341_ = branch_spec_i ? addr_i : _339_;
  assign instr_addr = valid_req_q ? stored_addr_q : _341_;
  assign rdata_outstanding_s = rvalid_or_pmp_err ? { 1'h0, rdata_outstanding_n[1] } : rdata_outstanding_n;
  assign branch_discard_s = rvalid_or_pmp_err ? { 1'h0, branch_discard_n[1] } : branch_discard_n;
  assign rdata_pmp_err_s = rvalid_or_pmp_err ? { 1'h0, rdata_pmp_err_n[1] } : rdata_pmp_err_n;
  assign fifo_addr = branch_i ? addr_i : 32'd0;
  paramodauxy_ibex_fetch_fifoNUM_REQS3200000000000000000000000000000010  fifo_i (
    .busy_o(fifo_busy),
    .busy_o_t0(fifo_busy_t0),
    .clear_i(branch_or_mispredict),
    .clear_i_t0(branch_or_mispredict_t0),
    .clk_i(clk_i),
    .in_addr_i(fifo_addr),
    .in_addr_i_t0(fifo_addr_t0),
    .in_err_i(instr_or_pmp_err),
    .in_err_i_t0(instr_or_pmp_err_t0),
    .in_rdata_i(instr_rdata_i),
    .in_rdata_i_t0(instr_rdata_i_t0),
    .in_valid_i(fifo_valid),
    .in_valid_i_t0(fifo_valid_t0),
    .out_addr_next_o(addr_next),
    .out_addr_next_o_t0(addr_next_t0),
    .out_addr_o(addr_o),
    .out_addr_o_t0(addr_o_t0),
    .out_err_o(err_o),
    .out_err_o_t0(err_o_t0),
    .out_err_plus2_o(err_plus2_o),
    .out_err_plus2_o_t0(err_plus2_o_t0),
    .out_rdata_o(rdata_o),
    .out_rdata_o_t0(rdata_o_t0),
    .out_ready_i(ready_i),
    .out_ready_i_t0(ready_i_t0),
    .out_valid_o(valid_raw),
    .out_valid_o_t0(valid_raw_t0),
    .rst_ni(rst_ni)
  );
  assign instr_addr_o = { instr_addr[31:2], 2'h0 };
  assign instr_addr_o_t0 = { instr_addr_t0[31:2], 2'h0 };
endmodule

module paramodauxy_ibex_wb_stageWritebackStage11 (clk_i, rst_ni, en_wb_i, instr_type_wb_i, pc_id_i, instr_is_compressed_id_i, instr_perf_count_id_i, ready_wb_o, rf_write_wb_o, outstanding_load_wb_o, outstanding_store_wb_o, pc_wb_o, perf_instr_ret_wb_o, perf_instr_ret_compressed_wb_o, rf_waddr_id_i, rf_wdata_id_i, rf_we_id_i, rf_wdata_lsu_i, rf_we_lsu_i, rf_wdata_fwd_wb_o, rf_waddr_wb_o
, rf_wdata_wb_o, rf_we_wb_o, lsu_resp_valid_i, lsu_resp_err_i, instr_done_wb_o, pc_id_i_t0, lsu_resp_valid_i_t0, en_wb_i_t0, instr_done_wb_o_t0, instr_is_compressed_id_i_t0, instr_perf_count_id_i_t0, instr_type_wb_i_t0, lsu_resp_err_i_t0, outstanding_load_wb_o_t0, outstanding_store_wb_o_t0, pc_wb_o_t0, perf_instr_ret_compressed_wb_o_t0, perf_instr_ret_wb_o_t0, ready_wb_o_t0, rf_waddr_id_i_t0, rf_waddr_wb_o_t0
, rf_wdata_fwd_wb_o_t0, rf_wdata_id_i_t0, rf_wdata_lsu_i_t0, rf_wdata_wb_o_t0, rf_we_id_i_t0, rf_we_lsu_i_t0, rf_we_wb_o_t0, rf_write_wb_o_t0);
  wire _000_;
  wire _001_;
  wire _002_;
  wire _003_;
  wire _004_;
  wire _005_;
  wire _006_;
  wire _007_;
  wire [1:0] _008_;
  wire _009_;
  wire _010_;
  wire _011_;
  wire _012_;
  wire _013_;
  wire _014_;
  wire _015_;
  wire [1:0] _016_;
  wire [31:0] _017_;
  wire _018_;
  wire _019_;
  wire _020_;
  wire _021_;
  wire _022_;
  wire _023_;
  wire _024_;
  wire _025_;
  wire _026_;
  wire _027_;
  wire _028_;
  wire _029_;
  wire _030_;
  wire _031_;
  wire _032_;
  wire _033_;
  wire _034_;
  wire _035_;
  wire _036_;
  wire _037_;
  wire _038_;
  wire _039_;
  wire _040_;
  wire _041_;
  wire _042_;
  wire _043_;
  wire _044_;
  wire _045_;
  wire _046_;
  wire _047_;
  wire _048_;
  wire _049_;
  wire _050_;
  wire _051_;
  wire _052_;
  wire [31:0] _053_;
  wire [31:0] _054_;
  wire [31:0] _055_;
  wire _056_;
  wire _057_;
  wire _058_;
  wire [4:0] _059_;
  wire [4:0] _060_;
  wire [4:0] _061_;
  wire [31:0] _062_;
  wire [31:0] _063_;
  wire [31:0] _064_;
  wire _065_;
  wire _066_;
  wire _067_;
  wire _068_;
  wire _069_;
  wire _070_;
  wire [1:0] _071_;
  wire [1:0] _072_;
  wire [1:0] _073_;
  wire [1:0] _074_;
  wire [1:0] _075_;
  wire [1:0] _076_;
  wire _077_;
  wire _078_;
  wire _079_;
  wire _080_;
  wire _081_;
  wire _082_;
  wire _083_;
  wire _084_;
  wire _085_;
  wire [1:0] _086_;
  wire [31:0] _087_;
  wire [31:0] _088_;
  wire [31:0] _089_;
  wire _090_;
  wire _091_;
  wire _092_;
  wire _093_;
  wire _094_;
  wire _095_;
  wire _096_;
  wire _097_;
  wire _098_;
  wire _099_;
  wire _100_;
  wire [31:0] _101_;
  wire [31:0] _102_;
  wire [31:0] _103_;
  wire [31:0] _104_;
  wire _105_;
  wire _106_;
  wire _107_;
  wire _108_;
  wire [4:0] _109_;
  wire [4:0] _110_;
  wire [4:0] _111_;
  wire [4:0] _112_;
  wire [31:0] _113_;
  wire [31:0] _114_;
  wire [31:0] _115_;
  wire [31:0] _116_;
  wire _117_;
  wire _118_;
  wire _119_;
  wire _120_;
  wire _121_;
  wire _122_;
  wire _123_;
  wire _124_;
  wire [1:0] _125_;
  wire [1:0] _126_;
  wire [1:0] _127_;
  wire [1:0] _128_;
  wire _129_;
  wire _130_;
  wire _131_;
  wire [31:0] _132_;
  wire [31:0] _133_;
  wire [31:0] _134_;
  wire [31:0] _135_;
  wire _136_;
  wire [4:0] _137_;
  wire [31:0] _138_;
  wire _139_;
  wire _140_;
  wire [1:0] _141_;
  wire [31:0] _142_;
  wire _143_;
  wire _144_;
  wire _145_;
  wire _146_;
  wire _147_;
  wire _148_;
  wire _149_;
  wire _150_;
  wire _151_;
  wire _152_;
  wire _153_;
  wire _154_;
  input clk_i;
  wire clk_i;
  input en_wb_i;
  wire en_wb_i;
  input en_wb_i_t0;
  wire en_wb_i_t0;
  reg \g_writeback_stage.rf_we_wb_q ;
  reg \g_writeback_stage.rf_we_wb_q_t0 ;
  reg \g_writeback_stage.wb_compressed_q ;
  reg \g_writeback_stage.wb_compressed_q_t0 ;
  reg \g_writeback_stage.wb_count_q ;
  reg \g_writeback_stage.wb_count_q_t0 ;
  wire \g_writeback_stage.wb_done ;
  wire \g_writeback_stage.wb_done_t0 ;
  reg [1:0] \g_writeback_stage.wb_instr_type_q ;
  reg [1:0] \g_writeback_stage.wb_instr_type_q_t0 ;
  wire \g_writeback_stage.wb_valid_d ;
  wire \g_writeback_stage.wb_valid_d_t0 ;
  reg \g_writeback_stage.wb_valid_q ;
  reg \g_writeback_stage.wb_valid_q_t0 ;
  output instr_done_wb_o;
  wire instr_done_wb_o;
  output instr_done_wb_o_t0;
  wire instr_done_wb_o_t0;
  input instr_is_compressed_id_i;
  wire instr_is_compressed_id_i;
  input instr_is_compressed_id_i_t0;
  wire instr_is_compressed_id_i_t0;
  input instr_perf_count_id_i;
  wire instr_perf_count_id_i;
  input instr_perf_count_id_i_t0;
  wire instr_perf_count_id_i_t0;
  input [1:0] instr_type_wb_i;
  wire [1:0] instr_type_wb_i;
  input [1:0] instr_type_wb_i_t0;
  wire [1:0] instr_type_wb_i_t0;
  input lsu_resp_err_i;
  wire lsu_resp_err_i;
  input lsu_resp_err_i_t0;
  wire lsu_resp_err_i_t0;
  input lsu_resp_valid_i;
  wire lsu_resp_valid_i;
  input lsu_resp_valid_i_t0;
  wire lsu_resp_valid_i_t0;
  output outstanding_load_wb_o;
  wire outstanding_load_wb_o;
  output outstanding_load_wb_o_t0;
  wire outstanding_load_wb_o_t0;
  output outstanding_store_wb_o;
  wire outstanding_store_wb_o;
  output outstanding_store_wb_o_t0;
  wire outstanding_store_wb_o_t0;
  input [31:0] pc_id_i;
  wire [31:0] pc_id_i;
  input [31:0] pc_id_i_t0;
  wire [31:0] pc_id_i_t0;
  output [31:0] pc_wb_o;
  reg [31:0] pc_wb_o;
  output [31:0] pc_wb_o_t0;
  reg [31:0] pc_wb_o_t0;
  output perf_instr_ret_compressed_wb_o;
  wire perf_instr_ret_compressed_wb_o;
  output perf_instr_ret_compressed_wb_o_t0;
  wire perf_instr_ret_compressed_wb_o_t0;
  output perf_instr_ret_wb_o;
  wire perf_instr_ret_wb_o;
  output perf_instr_ret_wb_o_t0;
  wire perf_instr_ret_wb_o_t0;
  output ready_wb_o;
  wire ready_wb_o;
  output ready_wb_o_t0;
  wire ready_wb_o_t0;
  input [4:0] rf_waddr_id_i;
  wire [4:0] rf_waddr_id_i;
  input [4:0] rf_waddr_id_i_t0;
  wire [4:0] rf_waddr_id_i_t0;
  output [4:0] rf_waddr_wb_o;
  reg [4:0] rf_waddr_wb_o;
  output [4:0] rf_waddr_wb_o_t0;
  reg [4:0] rf_waddr_wb_o_t0;
  output [31:0] rf_wdata_fwd_wb_o;
  reg [31:0] rf_wdata_fwd_wb_o;
  output [31:0] rf_wdata_fwd_wb_o_t0;
  reg [31:0] rf_wdata_fwd_wb_o_t0;
  input [31:0] rf_wdata_id_i;
  wire [31:0] rf_wdata_id_i;
  input [31:0] rf_wdata_id_i_t0;
  wire [31:0] rf_wdata_id_i_t0;
  input [31:0] rf_wdata_lsu_i;
  wire [31:0] rf_wdata_lsu_i;
  input [31:0] rf_wdata_lsu_i_t0;
  wire [31:0] rf_wdata_lsu_i_t0;
  wire [1:0] rf_wdata_wb_mux_we;
  wire [1:0] rf_wdata_wb_mux_we_t0;
  output [31:0] rf_wdata_wb_o;
  wire [31:0] rf_wdata_wb_o;
  output [31:0] rf_wdata_wb_o_t0;
  wire [31:0] rf_wdata_wb_o_t0;
  input rf_we_id_i;
  wire rf_we_id_i;
  input rf_we_id_i_t0;
  wire rf_we_id_i_t0;
  input rf_we_lsu_i;
  wire rf_we_lsu_i;
  input rf_we_lsu_i_t0;
  wire rf_we_lsu_i_t0;
  output rf_we_wb_o;
  wire rf_we_wb_o;
  output rf_we_wb_o_t0;
  wire rf_we_wb_o_t0;
  output rf_write_wb_o;
  wire rf_write_wb_o;
  output rf_write_wb_o_t0;
  wire rf_write_wb_o_t0;
  input rst_ni;
  wire rst_ni;
  assign _000_ = en_wb_i & ready_wb_o;
  assign _002_ = \g_writeback_stage.wb_valid_q  & _013_;
  assign rf_wdata_wb_mux_we[0] = \g_writeback_stage.rf_we_wb_q  & \g_writeback_stage.wb_valid_q ;
  assign rf_write_wb_o = \g_writeback_stage.wb_valid_q  & _153_;
  assign outstanding_load_wb_o = \g_writeback_stage.wb_valid_q  & _147_;
  assign outstanding_store_wb_o = \g_writeback_stage.wb_valid_q  & _149_;
  assign instr_done_wb_o = \g_writeback_stage.wb_valid_q  & \g_writeback_stage.wb_done ;
  assign _003_ = instr_done_wb_o & \g_writeback_stage.wb_count_q ;
  assign _005_ = lsu_resp_valid_i & lsu_resp_err_i;
  assign perf_instr_ret_wb_o = _003_ & _152_;
  assign perf_instr_ret_compressed_wb_o = perf_instr_ret_wb_o & \g_writeback_stage.wb_compressed_q ;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) \g_writeback_stage.wb_valid_q_t0  <= 1'h0;
    else \g_writeback_stage.wb_valid_q_t0  <= \g_writeback_stage.wb_valid_d_t0 ;
  assign _022_ = en_wb_i_t0 & ready_wb_o;
  assign _028_ = \g_writeback_stage.rf_we_wb_q_t0  & \g_writeback_stage.wb_valid_q ;
  assign _031_ = \g_writeback_stage.wb_valid_q_t0  & _153_;
  assign _034_ = \g_writeback_stage.wb_valid_q_t0  & _147_;
  assign _037_ = \g_writeback_stage.wb_valid_q_t0  & _149_;
  assign _040_ = \g_writeback_stage.wb_valid_q_t0  & \g_writeback_stage.wb_done ;
  assign _041_ = instr_done_wb_o_t0 & \g_writeback_stage.wb_count_q ;
  assign _044_ = lsu_resp_valid_i_t0 & lsu_resp_err_i;
  assign _047_ = _004_ & _152_;
  assign _050_ = perf_instr_ret_wb_o_t0 & \g_writeback_stage.wb_compressed_q ;
  assign _023_ = ready_wb_o_t0 & en_wb_i;
  assign _029_ = \g_writeback_stage.wb_valid_q_t0  & \g_writeback_stage.rf_we_wb_q ;
  assign _032_ = _154_ & \g_writeback_stage.wb_valid_q ;
  assign _035_ = _148_ & \g_writeback_stage.wb_valid_q ;
  assign _038_ = _150_ & \g_writeback_stage.wb_valid_q ;
  assign _042_ = \g_writeback_stage.wb_count_q_t0  & instr_done_wb_o;
  assign _045_ = lsu_resp_err_i_t0 & lsu_resp_valid_i;
  assign _048_ = _006_ & _003_;
  assign _051_ = \g_writeback_stage.wb_compressed_q_t0  & perf_instr_ret_wb_o;
  assign _024_ = en_wb_i_t0 & ready_wb_o_t0;
  assign _030_ = \g_writeback_stage.rf_we_wb_q_t0  & \g_writeback_stage.wb_valid_q_t0 ;
  assign _033_ = \g_writeback_stage.wb_valid_q_t0  & _154_;
  assign _036_ = \g_writeback_stage.wb_valid_q_t0  & _148_;
  assign _039_ = \g_writeback_stage.wb_valid_q_t0  & _150_;
  assign _043_ = instr_done_wb_o_t0 & \g_writeback_stage.wb_count_q_t0 ;
  assign _046_ = lsu_resp_valid_i_t0 & lsu_resp_err_i_t0;
  assign _049_ = _004_ & _006_;
  assign _052_ = perf_instr_ret_wb_o_t0 & \g_writeback_stage.wb_compressed_q_t0 ;
  assign _090_ = _022_ | _023_;
  assign _092_ = _028_ | _029_;
  assign _093_ = _031_ | _032_;
  assign _094_ = _034_ | _035_;
  assign _095_ = _037_ | _038_;
  assign _096_ = _040_ | _026_;
  assign _097_ = _041_ | _042_;
  assign _098_ = _044_ | _045_;
  assign _099_ = _047_ | _048_;
  assign _100_ = _050_ | _051_;
  assign _001_ = _090_ | _024_;
  assign rf_wdata_wb_mux_we_t0[0] = _092_ | _030_;
  assign rf_write_wb_o_t0 = _093_ | _033_;
  assign outstanding_load_wb_o_t0 = _094_ | _036_;
  assign outstanding_store_wb_o_t0 = _095_ | _039_;
  assign instr_done_wb_o_t0 = _096_ | _027_;
  assign _004_ = _097_ | _043_;
  assign _006_ = _098_ | _046_;
  assign perf_instr_ret_wb_o_t0 = _099_ | _049_;
  assign perf_instr_ret_compressed_wb_o_t0 = _100_ | _052_;
  assign _135_ = rf_wdata_id_i ^ rf_wdata_fwd_wb_o;
  assign _136_ = rf_we_id_i ^ \g_writeback_stage.rf_we_wb_q ;
  assign _137_ = rf_waddr_id_i ^ rf_waddr_wb_o;
  assign _138_ = pc_id_i ^ pc_wb_o;
  assign _139_ = instr_is_compressed_id_i ^ \g_writeback_stage.wb_compressed_q ;
  assign _140_ = instr_perf_count_id_i ^ \g_writeback_stage.wb_count_q ;
  assign _141_ = instr_type_wb_i ^ \g_writeback_stage.wb_instr_type_q ;
  assign _007_ = ~ en_wb_i;
  assign _101_ = rf_wdata_id_i_t0 | rf_wdata_fwd_wb_o_t0;
  assign _105_ = rf_we_id_i_t0 | \g_writeback_stage.rf_we_wb_q_t0 ;
  assign _109_ = rf_waddr_id_i_t0 | rf_waddr_wb_o_t0;
  assign _113_ = pc_id_i_t0 | pc_wb_o_t0;
  assign _117_ = instr_is_compressed_id_i_t0 | \g_writeback_stage.wb_compressed_q_t0 ;
  assign _121_ = instr_perf_count_id_i_t0 | \g_writeback_stage.wb_count_q_t0 ;
  assign _125_ = instr_type_wb_i_t0 | \g_writeback_stage.wb_instr_type_q_t0 ;
  assign _102_ = _135_ | _101_;
  assign _106_ = _136_ | _105_;
  assign _110_ = _137_ | _109_;
  assign _114_ = _138_ | _113_;
  assign _118_ = _139_ | _117_;
  assign _122_ = _140_ | _121_;
  assign _126_ = _141_ | _125_;
  assign _053_ = { en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i } & rf_wdata_id_i_t0;
  assign _056_ = en_wb_i & rf_we_id_i_t0;
  assign _059_ = { en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i } & rf_waddr_id_i_t0;
  assign _062_ = { en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i } & pc_id_i_t0;
  assign _065_ = en_wb_i & instr_is_compressed_id_i_t0;
  assign _068_ = en_wb_i & instr_perf_count_id_i_t0;
  assign _071_ = { en_wb_i, en_wb_i } & instr_type_wb_i_t0;
  assign _054_ = { _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_ } & rf_wdata_fwd_wb_o_t0;
  assign _057_ = _007_ & \g_writeback_stage.rf_we_wb_q_t0 ;
  assign _060_ = { _007_, _007_, _007_, _007_, _007_ } & rf_waddr_wb_o_t0;
  assign _063_ = { _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_ } & pc_wb_o_t0;
  assign _066_ = _007_ & \g_writeback_stage.wb_compressed_q_t0 ;
  assign _069_ = _007_ & \g_writeback_stage.wb_count_q_t0 ;
  assign _072_ = { _007_, _007_ } & \g_writeback_stage.wb_instr_type_q_t0 ;
  assign _055_ = _102_ & en_wb_i_t0;
  assign _058_ = _106_ & en_wb_i_t0;
  assign _061_ = _110_ & en_wb_i_t0;
  assign _064_ = _114_ & en_wb_i_t0;
  assign _067_ = _118_ & en_wb_i_t0;
  assign _070_ = _122_ & en_wb_i_t0;
  assign _073_ = _126_ & en_wb_i_t0;
  assign _103_ = _053_ | _054_;
  assign _107_ = _056_ | _057_;
  assign _111_ = _059_ | _060_;
  assign _115_ = _062_ | _063_;
  assign _119_ = _065_ | _066_;
  assign _123_ = _068_ | _069_;
  assign _127_ = _071_ | _072_;
  assign _104_ = _103_ | _055_;
  assign _108_ = _107_ | _058_;
  assign _112_ = _111_ | _061_;
  assign _116_ = _115_ | _064_;
  assign _120_ = _119_ | _067_;
  assign _124_ = _123_ | _070_;
  assign _128_ = _127_ | _073_;
  always_ff @(posedge clk_i)
    rf_wdata_fwd_wb_o_t0 <= _104_;
  always_ff @(posedge clk_i)
    \g_writeback_stage.rf_we_wb_q_t0  <= _108_;
  always_ff @(posedge clk_i)
    rf_waddr_wb_o_t0 <= _112_;
  always_ff @(posedge clk_i)
    pc_wb_o_t0 <= _116_;
  always_ff @(posedge clk_i)
    \g_writeback_stage.wb_compressed_q_t0  <= _120_;
  always_ff @(posedge clk_i)
    \g_writeback_stage.wb_count_q_t0  <= _124_;
  always_ff @(posedge clk_i)
    \g_writeback_stage.wb_instr_type_q_t0  <= _128_;
  assign _018_ = | \g_writeback_stage.wb_instr_type_q_t0 ;
  assign _008_ = ~ \g_writeback_stage.wb_instr_type_q_t0 ;
  assign _074_ = \g_writeback_stage.wb_instr_type_q  & _008_;
  assign _075_ = 2'h2 & _008_;
  assign _076_ = 2'h1 & _008_;
  assign _143_ = _074_ == _075_;
  assign _144_ = _074_ == _076_;
  assign _146_ = _143_ & _018_;
  assign _150_ = _144_ & _018_;
  always_ff @(posedge clk_i)
    if (en_wb_i) rf_wdata_fwd_wb_o <= rf_wdata_id_i;
  always_ff @(posedge clk_i)
    if (en_wb_i) \g_writeback_stage.rf_we_wb_q  <= rf_we_id_i;
  always_ff @(posedge clk_i)
    if (en_wb_i) rf_waddr_wb_o <= rf_waddr_id_i;
  always_ff @(posedge clk_i)
    if (en_wb_i) pc_wb_o <= pc_id_i;
  always_ff @(posedge clk_i)
    if (en_wb_i) \g_writeback_stage.wb_compressed_q  <= instr_is_compressed_id_i;
  always_ff @(posedge clk_i)
    if (en_wb_i) \g_writeback_stage.wb_count_q  <= instr_perf_count_id_i;
  always_ff @(posedge clk_i)
    if (en_wb_i) \g_writeback_stage.wb_instr_type_q  <= instr_type_wb_i;
  assign _019_ = | { rf_wdata_wb_mux_we_t0[0], rf_we_lsu_i_t0 };
  assign _016_ = ~ { rf_wdata_wb_mux_we_t0[0], rf_we_lsu_i_t0 };
  assign _086_ = { rf_wdata_wb_mux_we[0], rf_we_lsu_i } & _016_;
  assign _020_ = ! _074_;
  assign _021_ = ! _086_;
  assign _148_ = _020_ & _018_;
  assign rf_we_wb_o_t0 = _021_ & _019_;
  assign _017_ = ~ { rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0] };
  assign _132_ = { rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0] } | _017_;
  assign _133_ = { rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0] } | { rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0] };
  assign _087_ = rf_wdata_lsu_i_t0 & _132_;
  assign _088_ = rf_wdata_fwd_wb_o_t0 & _133_;
  assign _134_ = _087_ | _088_;
  assign _142_ = rf_wdata_lsu_i ^ rf_wdata_fwd_wb_o;
  assign _089_ = { rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0] } & _142_;
  assign rf_wdata_wb_o_t0 = _089_ | _134_;
  assign _009_ = ~ _000_;
  assign _011_ = ~ _145_;
  assign _014_ = ~ \g_writeback_stage.rf_we_wb_q ;
  assign _010_ = ~ _002_;
  assign _012_ = ~ lsu_resp_valid_i;
  assign _013_ = ~ \g_writeback_stage.wb_done ;
  assign _015_ = ~ _147_;
  assign _077_ = _001_ & _010_;
  assign _080_ = _146_ & _012_;
  assign _025_ = \g_writeback_stage.wb_valid_q_t0  & _013_;
  assign _083_ = \g_writeback_stage.rf_we_wb_q_t0  & _015_;
  assign _078_ = ready_wb_o_t0 & _009_;
  assign _081_ = lsu_resp_valid_i_t0 & _011_;
  assign _026_ = \g_writeback_stage.wb_done_t0  & \g_writeback_stage.wb_valid_q ;
  assign _084_ = _148_ & _014_;
  assign _079_ = _001_ & ready_wb_o_t0;
  assign _082_ = _146_ & lsu_resp_valid_i_t0;
  assign _027_ = \g_writeback_stage.wb_valid_q_t0  & \g_writeback_stage.wb_done_t0 ;
  assign _085_ = \g_writeback_stage.rf_we_wb_q_t0  & _148_;
  assign _129_ = _077_ | _078_;
  assign _130_ = _080_ | _081_;
  assign _091_ = _025_ | _026_;
  assign _131_ = _083_ | _084_;
  assign \g_writeback_stage.wb_valid_d_t0  = _129_ | _079_;
  assign \g_writeback_stage.wb_done_t0  = _130_ | _082_;
  assign ready_wb_o_t0 = _091_ | _027_;
  assign _154_ = _131_ | _085_;
  assign _145_ = \g_writeback_stage.wb_instr_type_q  == 2'h2;
  assign _147_ = ! \g_writeback_stage.wb_instr_type_q ;
  assign _149_ = \g_writeback_stage.wb_instr_type_q  == 2'h1;
  assign _151_ = ~ \g_writeback_stage.wb_valid_q ;
  assign _152_ = ~ _005_;
  assign \g_writeback_stage.wb_valid_d  = _000_ | _002_;
  assign \g_writeback_stage.wb_done  = _145_ | lsu_resp_valid_i;
  assign ready_wb_o = _151_ | \g_writeback_stage.wb_done ;
  assign _153_ = \g_writeback_stage.rf_we_wb_q  | _147_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) \g_writeback_stage.wb_valid_q  <= 1'h0;
    else \g_writeback_stage.wb_valid_q  <= \g_writeback_stage.wb_valid_d ;
  assign rf_we_wb_o = | { rf_wdata_wb_mux_we[0], rf_we_lsu_i };
  assign rf_wdata_wb_o = rf_wdata_wb_mux_we[0] ? rf_wdata_fwd_wb_o : rf_wdata_lsu_i;
  assign rf_wdata_wb_mux_we[1] = rf_we_lsu_i;
  assign rf_wdata_wb_mux_we_t0[1] = rf_we_lsu_i_t0;
endmodule

module paramodauxy_prim_diff_decodeAsyncOn10 (clk_i, rst_ni, diff_pi, diff_ni, level_o, rise_o, fall_o, event_o, sigint_o, diff_ni_t0, diff_pi_t0, event_o_t0, fall_o_t0, level_o_t0, rise_o_t0, sigint_o_t0);
  wire _00_;
  wire _01_;
  wire _02_;
  wire _03_;
  wire _04_;
  wire _05_;
  wire _06_;
  wire _07_;
  wire _08_;
  wire _09_;
  wire _10_;
  wire _11_;
  wire _12_;
  wire _13_;
  wire _14_;
  wire _15_;
  wire _16_;
  wire _17_;
  wire _18_;
  wire _19_;
  wire _20_;
  wire _21_;
  wire _22_;
  wire _23_;
  wire _24_;
  wire _25_;
  wire _26_;
  wire _27_;
  wire _28_;
  wire _29_;
  wire _30_;
  wire _31_;
  wire _32_;
  wire _33_;
  wire _34_;
  input clk_i;
  wire clk_i;
  input diff_ni;
  wire diff_ni;
  input diff_ni_t0;
  wire diff_ni_t0;
  input diff_pi;
  wire diff_pi;
  input diff_pi_t0;
  wire diff_pi_t0;
  output event_o;
  wire event_o;
  output event_o_t0;
  wire event_o_t0;
  output fall_o;
  wire fall_o;
  output fall_o_t0;
  wire fall_o_t0;
  reg \gen_no_async.diff_pq ;
  reg \gen_no_async.diff_pq_t0 ;
  output level_o;
  wire level_o;
  output level_o_t0;
  wire level_o_t0;
  reg level_q;
  reg level_q_t0;
  output rise_o;
  wire rise_o;
  output rise_o_t0;
  wire rise_o_t0;
  input rst_ni;
  wire rst_ni;
  output sigint_o;
  wire sigint_o;
  output sigint_o_t0;
  wire sigint_o_t0;
  assign _00_ = _32_ & diff_pi;
  assign rise_o = _00_ & _33_;
  assign _02_ = \gen_no_async.diff_pq  & _34_;
  assign fall_o = _02_ & _33_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) level_q_t0 <= 1'h0;
    else level_q_t0 <= level_o_t0;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) \gen_no_async.diff_pq_t0  <= 1'h0;
    else \gen_no_async.diff_pq_t0  <= diff_pi_t0;
  assign _06_ = \gen_no_async.diff_pq_t0  & diff_pi;
  assign _09_ = _01_ & _33_;
  assign _12_ = \gen_no_async.diff_pq_t0  & _34_;
  assign _14_ = _03_ & _33_;
  assign _07_ = diff_pi_t0 & _32_;
  assign _10_ = sigint_o_t0 & _00_;
  assign _13_ = diff_pi_t0 & \gen_no_async.diff_pq ;
  assign _15_ = sigint_o_t0 & _02_;
  assign _11_ = _01_ & sigint_o_t0;
  assign _08_ = \gen_no_async.diff_pq_t0  & diff_pi_t0;
  assign _16_ = _03_ & sigint_o_t0;
  assign _23_ = _06_ | _07_;
  assign _24_ = _09_ | _10_;
  assign _25_ = _12_ | _13_;
  assign _26_ = _14_ | _15_;
  assign _01_ = _23_ | _08_;
  assign rise_o_t0 = _24_ | _11_;
  assign _03_ = _25_ | _08_;
  assign fall_o_t0 = _26_ | _16_;
  assign sigint_o = ~ _33_;
  assign _28_ = sigint_o_t0 | sigint_o;
  assign _29_ = sigint_o_t0 | _33_;
  assign _20_ = level_q_t0 & _28_;
  assign _21_ = diff_pi_t0 & _29_;
  assign _30_ = _20_ | _21_;
  assign _31_ = level_q ^ diff_pi;
  assign _22_ = sigint_o_t0 & _31_;
  assign level_o_t0 = _22_ | _30_;
  assign _04_ = ~ rise_o;
  assign _05_ = ~ fall_o;
  assign _17_ = rise_o_t0 & _05_;
  assign _18_ = fall_o_t0 & _04_;
  assign _19_ = rise_o_t0 & fall_o_t0;
  assign _27_ = _17_ | _18_;
  assign event_o_t0 = _27_ | _19_;
  assign sigint_o_t0 = diff_pi_t0 | diff_ni_t0;
  assign _32_ = ~ \gen_no_async.diff_pq ;
  assign _34_ = ~ diff_pi;
  assign event_o = rise_o | fall_o;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) level_q <= 1'h0;
    else level_q <= level_o;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) \gen_no_async.diff_pq  <= 1'h0;
    else \gen_no_async.diff_pq  <= diff_pi;
  assign level_o = _33_ ? diff_pi : level_q;
  assign _33_ = diff_pi ^ diff_ni;
endmodule





module paramodauxy_prim_flopWidths3200000000000000000000000000000001ResetValue10 (clk_i, rst_ni, d_i, q_o, q_o_t0, d_i_t0);
  input clk_i;
  wire clk_i;
  input d_i;
  wire d_i;
  input d_i_t0;
  wire d_i_t0;
  output q_o;
  wire q_o;
  output q_o_t0;
  wire q_o_t0;
  input rst_ni;
  wire rst_ni;
  paramodauxy_prim_generic_flopWidths3200000000000000000000000000000001ResetValue10  \gen_generic.u_impl_generic  (
    .clk_i(clk_i),
    .d_i(d_i),
    .d_i_t0(d_i_t0),
    .q_o(q_o),
    .q_o_t0(q_o_t0),
    .rst_ni(rst_ni)
  );
endmodule

module paramodauxy_prim_flop_2syncWidths3200000000000000000000000000000001 (clk_i, rst_ni, d_i, q_o, q_o_t0, d_i_t0);
  input clk_i;
  wire clk_i;
  input d_i;
  wire d_i;
  input d_i_t0;
  wire d_i_t0;
  output q_o;
  wire q_o;
  output q_o_t0;
  wire q_o_t0;
  input rst_ni;
  wire rst_ni;
  paramodauxy_prim_generic_flop_2syncWidths3200000000000000000000000000000001ResetValue10  \gen_generic.u_impl_generic  (
    .clk_i(clk_i),
    .d_i(d_i),
    .d_i_t0(d_i_t0),
    .q_o(q_o),
    .q_o_t0(q_o_t0),
    .rst_ni(rst_ni)
  );
endmodule

module paramodauxy_prim_generic_bufWidths3200000000000000000000000000000001 (in_i, out_o, in_i_t0, out_o_t0);
  input in_i;
  wire in_i;
  input in_i_t0;
  wire in_i_t0;
  output out_o;
  wire out_o;
  output out_o_t0;
  wire out_o_t0;
  assign out_o = in_i;
  assign out_o_t0 = in_i_t0;
endmodule

module paramodauxy_prim_generic_flopWidths3200000000000000000000000000000001ResetValue10 (clk_i, rst_ni, d_i, q_o, q_o_t0, d_i_t0);
  input clk_i;
  wire clk_i;
  input d_i;
  wire d_i;
  input d_i_t0;
  wire d_i_t0;
  output q_o;
  reg q_o;
  output q_o_t0;
  reg q_o_t0;
  input rst_ni;
  wire rst_ni;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) q_o_t0 <= 1'h0;
    else q_o_t0 <= d_i_t0;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) q_o <= 1'h0;
    else q_o <= d_i;
endmodule

module paramodauxy_prim_generic_flop_2syncWidths3200000000000000000000000000000001ResetValue10 (clk_i, rst_ni, d_i, q_o, q_o_t0, d_i_t0);
  input clk_i;
  wire clk_i;
  input d_i;
  wire d_i;
  input d_i_t0;
  wire d_i_t0;
  wire intq;
  wire intq_t0;
  output q_o;
  wire q_o;
  output q_o_t0;
  wire q_o_t0;
  input rst_ni;
  wire rst_ni;
  paramodauxy_prim_flopWidths3200000000000000000000000000000001ResetValue10  u_sync_1 (
    .clk_i(clk_i),
    .d_i(d_i),
    .d_i_t0(d_i_t0),
    .q_o(intq),
    .q_o_t0(intq_t0),
    .rst_ni(rst_ni)
  );
  paramodauxy_prim_flopWidths3200000000000000000000000000000001ResetValue10  u_sync_2 (
    .clk_i(clk_i),
    .d_i(intq),
    .d_i_t0(intq_t0),
    .q_o(q_o),
    .q_o_t0(q_o_t0),
    .rst_ni(rst_ni)
  );
endmodule

module paramodauxy_tlul_adapter_hostMAX_REQSs3200000000000000000000000000000010 (clk_i, rst_ni, req_i, gnt_o, addr_i, we_i, wdata_i, be_i, type_i, valid_o, rdata_o, err_o, intg_err_o, tl_o, tl_i, wdata_i_t0, valid_o_t0, req_i_t0, err_o_t0, addr_i_t0, rdata_o_t0
, tl_i_t0, tl_o_t0, be_i_t0, gnt_o_t0, intg_err_o_t0, type_i_t0, we_i_t0);
  wire _000_;
  wire _001_;
  wire [31:0] _002_;
  wire [31:0] _003_;
  wire [31:0] _004_;
  wire _005_;
  wire _006_;
  wire _007_;
  wire _008_;
  wire _009_;
  wire [3:0] _010_;
  wire [2:0] _011_;
  wire [2:0] _012_;
  wire _013_;
  wire _014_;
  wire [31:0] _015_;
  wire _016_;
  wire _017_;
  wire _018_;
  wire _019_;
  wire _020_;
  wire _021_;
  wire _022_;
  wire _023_;
  wire _024_;
  wire _025_;
  wire _026_;
  wire _027_;
  wire _028_;
  wire _029_;
  wire _030_;
  wire [3:0] _031_;
  wire [3:0] _032_;
  wire [3:0] _033_;
  wire [2:0] _034_;
  wire [2:0] _035_;
  wire [2:0] _036_;
  wire [2:0] _037_;
  wire [2:0] _038_;
  wire [2:0] _039_;
  wire [31:0] _040_;
  wire _041_;
  wire _042_;
  wire _043_;
  wire _044_;
  wire _045_;
  wire _046_;
  wire _047_;
  wire _048_;
  wire _049_;
  wire _050_;
  wire [3:0] _051_;
  wire [3:0] _052_;
  wire [3:0] _053_;
  wire [3:0] _054_;
  wire [2:0] _055_;
  wire [2:0] _056_;
  wire [2:0] _057_;
  wire [2:0] _058_;
  wire [2:0] _059_;
  wire [2:0] _060_;
  wire [31:0] _061_;
  wire _062_;
  wire [3:0] _063_;
  wire [2:0] _064_;
  wire [31:0] _065_;
  wire [31:0] _066_;
  wire _067_;
  wire _068_;
  wire _069_;
  wire _070_;
  wire [2:0] _071_;
  wire [2:0] _072_;
  input [31:0] addr_i;
  wire [31:0] addr_i;
  input [31:0] addr_i_t0;
  wire [31:0] addr_i_t0;
  input [3:0] be_i;
  wire [3:0] be_i;
  input [3:0] be_i_t0;
  wire [3:0] be_i_t0;
  input clk_i;
  wire clk_i;
  output err_o;
  wire err_o;
  output err_o_t0;
  wire err_o_t0;
  reg \g_multiple_reqs.source_q ;
  reg \g_multiple_reqs.source_q_t0 ;
  output gnt_o;
  wire gnt_o;
  output gnt_o_t0;
  wire gnt_o_t0;
  wire intg_err;
  output intg_err_o;
  wire intg_err_o;
  output intg_err_o_t0;
  wire intg_err_o_t0;
  reg intg_err_q;
  reg intg_err_q_t0;
  wire intg_err_t0;
  output [31:0] rdata_o;
  wire [31:0] rdata_o;
  output [31:0] rdata_o_t0;
  wire [31:0] rdata_o_t0;
  input req_i;
  wire req_i;
  input req_i_t0;
  wire req_i_t0;
  input rst_ni;
  wire rst_ni;
  wire [3:0] tl_be;
  wire [3:0] tl_be_t0;
  input [65:0] tl_i;
  wire [65:0] tl_i;
  input [65:0] tl_i_t0;
  wire [65:0] tl_i_t0;
  output [106:0] tl_o;
  wire [106:0] tl_o;
  output [106:0] tl_o_t0;
  wire [106:0] tl_o_t0;
  wire [106:0] tl_out;
  wire [106:0] tl_out_t0;
  input [1:0] type_i;
  wire [1:0] type_i;
  input [1:0] type_i_t0;
  wire [1:0] type_i_t0;
  output valid_o;
  wire valid_o;
  output valid_o_t0;
  wire valid_o_t0;
  input [31:0] wdata_i;
  wire [31:0] wdata_i;
  input [31:0] wdata_i_t0;
  wire [31:0] wdata_i_t0;
  input we_i;
  wire we_i;
  input we_i_t0;
  wire we_i_t0;
  assign _002_ = \g_multiple_reqs.source_q  + 32'd1;
  assign _004_ = ~ { 31'h00000000, \g_multiple_reqs.source_q_t0  };
  assign _015_ = { 31'h00000000, \g_multiple_reqs.source_q  } & _004_;
  assign _065_ = _015_ + 32'd1;
  assign _040_ = { 31'h00000000, \g_multiple_reqs.source_q  } | { 31'h00000000, \g_multiple_reqs.source_q_t0  };
  assign _066_ = _040_ + 32'd1;
  assign _061_ = _065_ ^ _066_;
  assign _003_ = _061_ | { 31'h00000000, \g_multiple_reqs.source_q_t0  };
  assign _005_ = ~ _067_;
  assign _062_ = _000_ ^ \g_multiple_reqs.source_q ;
  assign _041_ = _001_ | \g_multiple_reqs.source_q_t0 ;
  assign _042_ = _062_ | _041_;
  assign _045_ = _008_ | intg_err_q_t0;
  assign _016_ = _067_ & _001_;
  assign _017_ = _005_ & \g_multiple_reqs.source_q_t0 ;
  assign _018_ = _042_ & _068_;
  assign _020_ = _045_ & intg_err_t0;
  assign _043_ = _016_ | _017_;
  assign _044_ = _043_ | _018_;
  assign _046_ = _019_ | _020_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) \g_multiple_reqs.source_q_t0  <= 1'h0;
    else \g_multiple_reqs.source_q_t0  <= _044_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) intg_err_q_t0 <= 1'h0;
    else intg_err_q_t0 <= _046_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) \g_multiple_reqs.source_q  <= 1'h0;
    else if (_067_) \g_multiple_reqs.source_q  <= _000_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) intg_err_q <= 1'h0;
    else if (intg_err) intg_err_q <= 1'h1;
  assign _021_ = req_i_t0 & tl_i[0];
  assign _022_ = tl_i_t0[0] & req_i;
  assign _023_ = req_i_t0 & tl_i_t0[0];
  assign _047_ = _021_ | _022_;
  assign _068_ = _047_ | _023_;
  assign _009_ = ~ \g_multiple_reqs.source_q ;
  assign _010_ = ~ { we_i, we_i, we_i, we_i };
  assign _011_ = ~ { _069_, _069_, _069_ };
  assign _012_ = ~ { we_i, we_i, we_i };
  assign _050_ = \g_multiple_reqs.source_q_t0  | _009_;
  assign _052_ = { we_i_t0, we_i_t0, we_i_t0, we_i_t0 } | _010_;
  assign _055_ = { _070_, _070_, _070_ } | _011_;
  assign _058_ = { we_i_t0, we_i_t0, we_i_t0 } | _012_;
  assign _053_ = { we_i_t0, we_i_t0, we_i_t0, we_i_t0 } | { we_i, we_i, we_i, we_i };
  assign _056_ = { _070_, _070_, _070_ } | { _069_, _069_, _069_ };
  assign _059_ = { we_i_t0, we_i_t0, we_i_t0 } | { we_i, we_i, we_i };
  assign _029_ = _003_[0] & _050_;
  assign _031_ = 4'h0 & _052_;
  assign _034_ = 3'h0 & _055_;
  assign _037_ = 3'h0 & _058_;
  assign _032_ = be_i_t0 & _053_;
  assign _035_ = 3'h0 & _056_;
  assign _038_ = _072_ & _059_;
  assign _054_ = _031_ | _032_;
  assign _057_ = _034_ | _035_;
  assign _060_ = _037_ | _038_;
  assign _063_ = 4'hf ^ be_i;
  assign _064_ = 3'h4 ^ _071_;
  assign _030_ = \g_multiple_reqs.source_q_t0  & _002_[0];
  assign _033_ = { we_i_t0, we_i_t0, we_i_t0, we_i_t0 } & _063_;
  assign _036_ = { _070_, _070_, _070_ } & 3'h1;
  assign _039_ = { we_i_t0, we_i_t0, we_i_t0 } & _064_;
  assign _001_ = _030_ | _029_;
  assign tl_be_t0 = _033_ | _054_;
  assign _072_ = _036_ | _057_;
  assign tl_out_t0[105:103] = _039_ | _060_;
  assign _007_ = ~ tl_i[1];
  assign _008_ = ~ intg_err_q;
  assign _006_ = ~ intg_err;
  assign _024_ = tl_i_t0[1] & _006_;
  assign _019_ = intg_err_q_t0 & _006_;
  assign _025_ = intg_err_t0 & _007_;
  assign _027_ = intg_err_t0 & _008_;
  assign _026_ = tl_i_t0[1] & intg_err_t0;
  assign _028_ = intg_err_q_t0 & intg_err_t0;
  assign _048_ = _024_ | _025_;
  assign _049_ = _019_ | _027_;
  assign err_o_t0 = _048_ | _026_;
  assign intg_err_o_t0 = _049_ | _028_;
  assign _014_ = | be_i_t0;
  assign _051_ = be_i | be_i_t0;
  assign _013_ = & _051_;
  assign _070_ = _014_ & _013_;
  assign _067_ = req_i && tl_i[0];
  assign err_o = tl_i[1] | intg_err;
  assign intg_err_o = intg_err_q | intg_err;
  assign _000_ = \g_multiple_reqs.source_q  ? 1'h0 : _002_[0];
  assign _069_ = & be_i;
  assign tl_be = we_i ? be_i : 4'hf;
  assign _071_ = _069_ ? 3'h0 : 3'h1;
  assign tl_out[105:103] = we_i ? _071_ : 3'h4;
  auxy_tlul_cmd_intg_gen u_cmd_intg_gen (
    .tl_i({ req_i, tl_out[105:103], 12'h100, \g_multiple_reqs.source_q , addr_i[31:2], 2'h0, tl_be, wdata_i, 5'h00, type_i, 15'h0001 }),
    .tl_i_t0({ req_i_t0, tl_out_t0[105:103], 12'h000, \g_multiple_reqs.source_q_t0 , addr_i_t0[31:2], 2'h0, tl_be_t0, wdata_i_t0, 5'h00, type_i_t0, 15'h0000 }),
    .tl_o(tl_o),
    .tl_o_t0(tl_o_t0)
  );
  auxy_tlul_rsp_intg_chk u_rsp_chk (
    .err_o(intg_err),
    .err_o_t0(intg_err_t0),
    .tl_i(tl_i),
    .tl_i_t0(tl_i_t0)
  );
  assign gnt_o = tl_i[0];
  assign gnt_o_t0 = tl_i_t0[0];
  assign rdata_o = tl_i[47:16];
  assign rdata_o_t0 = tl_i_t0[47:16];
  assign { tl_out[106], tl_out[102:0] } = { req_i, 12'h100, \g_multiple_reqs.source_q , addr_i[31:2], 2'h0, tl_be, wdata_i, 5'h00, type_i, 15'h0001 };
  assign { tl_out_t0[106], tl_out_t0[102:0] } = { req_i_t0, 12'h000, \g_multiple_reqs.source_q_t0 , addr_i_t0[31:2], 2'h0, tl_be_t0, wdata_i_t0, 5'h00, type_i_t0, 15'h0000 };
  assign valid_o = tl_i[65];
  assign valid_o_t0 = tl_i_t0[65];
endmodule

module paramodauxy_tlul_rsp_intg_genEnableRspIntgGen10EnableDataIntgGen10 (tl_i, tl_o, tl_i_t0, tl_o_t0);
  input [65:0] tl_i;
  wire [65:0] tl_i;
  input [65:0] tl_i_t0;
  wire [65:0] tl_i_t0;
  output [65:0] tl_o;
  wire [65:0] tl_o;
  output [65:0] tl_o_t0;
  wire [65:0] tl_o_t0;
  assign tl_o = tl_i;
  assign tl_o_t0 = tl_i_t0;
endmodule

module auxy_ibex_compressed_decoder(clk_i, rst_ni, valid_i, instr_i, instr_o, is_compressed_o, illegal_instr_o, valid_i_t0, is_compressed_o_t0, instr_o_t0, instr_i_t0, illegal_instr_o_t0);
  wire _0000_;
  wire [31:0] _0001_;
  wire [31:0] _0002_;
  wire _0003_;
  wire _0004_;
  wire [31:0] _0005_;
  wire [31:0] _0006_;
  wire _0007_;
  wire _0008_;
  wire _0009_;
  wire _0010_;
  wire _0011_;
  wire _0012_;
  wire [31:0] _0013_;
  wire [31:0] _0014_;
  wire _0015_;
  wire _0016_;
  wire [31:0] _0017_;
  wire [31:0] _0018_;
  wire _0019_;
  wire _0020_;
  wire [31:0] _0021_;
  wire [31:0] _0022_;
  wire _0023_;
  wire _0024_;
  wire [31:0] _0025_;
  wire [31:0] _0026_;
  wire _0027_;
  wire _0028_;
  wire [31:0] _0029_;
  wire [31:0] _0030_;
  wire [31:0] _0031_;
  wire [31:0] _0032_;
  wire _0033_;
  wire _0034_;
  wire [31:0] _0035_;
  wire [31:0] _0036_;
  wire _0037_;
  wire _0038_;
  wire [31:0] _0039_;
  wire [31:0] _0040_;
  wire _0041_;
  wire _0042_;
  wire _0043_;
  wire _0044_;
  wire [1:0] _0045_;
  wire [5:0] _0046_;
  wire _0047_;
  wire _0048_;
  wire _0049_;
  wire _0050_;
  wire _0051_;
  wire _0052_;
  wire _0053_;
  wire [3:0] _0054_;
  wire _0055_;
  wire _0056_;
  wire _0057_;
  wire [31:0] _0058_;
  wire [31:0] _0059_;
  wire [31:0] _0060_;
  wire [31:0] _0061_;
  wire [31:0] _0062_;
  wire [31:0] _0063_;
  wire [31:0] _0064_;
  wire [31:0] _0065_;
  wire _0066_;
  wire _0067_;
  wire [31:0] _0068_;
  wire [31:0] _0069_;
  wire [31:0] _0070_;
  wire [31:0] _0071_;
  wire [31:0] _0072_;
  wire _0073_;
  wire _0074_;
  wire [31:0] _0075_;
  wire [31:0] _0076_;
  wire _0077_;
  wire _0078_;
  wire [31:0] _0079_;
  wire [31:0] _0080_;
  wire [31:0] _0081_;
  wire [7:0] _0082_;
  wire [4:0] _0083_;
  wire [5:0] _0084_;
  wire [4:0] _0085_;
  wire [1:0] _0086_;
  wire [31:0] _0087_;
  wire [31:0] _0088_;
  wire _0089_;
  wire _0090_;
  wire [31:0] _0091_;
  wire [3:0] _0092_;
  wire [3:0] _0093_;
  wire [2:0] _0094_;
  wire [1:0] _0095_;
  wire [31:0] _0096_;
  wire [1:0] _0097_;
  wire [1:0] _0098_;
  wire [4:0] _0099_;
  wire [2:0] _0100_;
  wire _0101_;
  wire _0102_;
  wire _0103_;
  wire _0104_;
  wire _0105_;
  wire _0106_;
  wire _0107_;
  wire _0108_;
  wire _0109_;
  wire _0110_;
  wire _0111_;
  wire _0112_;
  wire _0113_;
  wire _0114_;
  wire _0115_;
  wire _0116_;
  wire _0117_;
  wire _0118_;
  wire _0119_;
  wire _0120_;
  wire _0121_;
  wire _0122_;
  wire _0123_;
  wire _0124_;
  wire _0125_;
  wire _0126_;
  wire _0127_;
  wire _0128_;
  wire _0129_;
  wire _0130_;
  wire _0131_;
  wire _0132_;
  wire [1:0] _0133_;
  wire [5:0] _0134_;
  wire _0135_;
  wire _0136_;
  wire _0137_;
  wire _0138_;
  wire _0139_;
  wire _0140_;
  wire _0141_;
  wire _0142_;
  wire _0143_;
  wire _0144_;
  wire _0145_;
  wire _0146_;
  wire [3:0] _0147_;
  wire _0148_;
  wire _0149_;
  wire _0150_;
  wire _0151_;
  wire _0152_;
  wire _0153_;
  wire _0154_;
  wire _0155_;
  wire _0156_;
  wire _0157_;
  wire [31:0] _0158_;
  wire [31:0] _0159_;
  wire [31:0] _0160_;
  wire [31:0] _0161_;
  wire [31:0] _0162_;
  wire [31:0] _0163_;
  wire [31:0] _0164_;
  wire [31:0] _0165_;
  wire [31:0] _0166_;
  wire [31:0] _0167_;
  wire [31:0] _0168_;
  wire [31:0] _0169_;
  wire [31:0] _0170_;
  wire [31:0] _0171_;
  wire [31:0] _0172_;
  wire [31:0] _0173_;
  wire [31:0] _0174_;
  wire [31:0] _0175_;
  wire [31:0] _0176_;
  wire [31:0] _0177_;
  wire [31:0] _0178_;
  wire [31:0] _0179_;
  wire [31:0] _0180_;
  wire [31:0] _0181_;
  wire _0182_;
  wire _0183_;
  wire _0184_;
  wire _0185_;
  wire _0186_;
  wire [31:0] _0187_;
  wire [31:0] _0188_;
  wire [31:0] _0189_;
  wire [31:0] _0190_;
  wire [31:0] _0191_;
  wire [31:0] _0192_;
  wire [31:0] _0193_;
  wire [31:0] _0194_;
  wire [31:0] _0195_;
  wire [31:0] _0196_;
  wire [31:0] _0197_;
  wire [31:0] _0198_;
  wire [31:0] _0199_;
  wire [31:0] _0200_;
  wire [31:0] _0201_;
  wire [31:0] _0202_;
  wire [31:0] _0203_;
  wire [31:0] _0204_;
  wire [31:0] _0205_;
  wire [31:0] _0206_;
  wire [31:0] _0207_;
  wire _0208_;
  wire _0209_;
  wire _0210_;
  wire _0211_;
  wire _0212_;
  wire _0213_;
  wire _0214_;
  wire _0215_;
  wire _0216_;
  wire [31:0] _0217_;
  wire [31:0] _0218_;
  wire [31:0] _0219_;
  wire [31:0] _0220_;
  wire [31:0] _0221_;
  wire [31:0] _0222_;
  wire [31:0] _0223_;
  wire [31:0] _0224_;
  wire [31:0] _0225_;
  wire _0226_;
  wire _0227_;
  wire _0228_;
  wire _0229_;
  wire _0230_;
  wire _0231_;
  wire _0232_;
  wire _0233_;
  wire [31:0] _0234_;
  wire [31:0] _0235_;
  wire [31:0] _0236_;
  wire [31:0] _0237_;
  wire [31:0] _0238_;
  wire [31:0] _0239_;
  wire [31:0] _0240_;
  wire [31:0] _0241_;
  wire [31:0] _0242_;
  wire [7:0] _0243_;
  wire [4:0] _0244_;
  wire [4:0] _0245_;
  wire [5:0] _0246_;
  wire [4:0] _0247_;
  wire [1:0] _0248_;
  wire [1:0] _0249_;
  wire [31:0] _0250_;
  wire [31:0] _0251_;
  wire [31:0] _0252_;
  wire [31:0] _0253_;
  wire [31:0] _0254_;
  wire [31:0] _0255_;
  wire [31:0] _0256_;
  wire [31:0] _0257_;
  wire [31:0] _0258_;
  wire _0259_;
  wire _0260_;
  wire _0261_;
  wire _0262_;
  wire [31:0] _0263_;
  wire [31:0] _0264_;
  wire [31:0] _0265_;
  wire [3:0] _0266_;
  wire [3:0] _0267_;
  wire [2:0] _0268_;
  wire [2:0] _0269_;
  wire [2:0] _0270_;
  wire [2:0] _0271_;
  wire [2:0] _0272_;
  wire [2:0] _0273_;
  wire [2:0] _0274_;
  wire [2:0] _0275_;
  wire [1:0] _0276_;
  wire [1:0] _0277_;
  wire [1:0] _0278_;
  wire [31:0] _0279_;
  wire [31:0] _0280_;
  wire [31:0] _0281_;
  wire [1:0] _0282_;
  wire [1:0] _0283_;
  wire [4:0] _0284_;
  wire [2:0] _0285_;
  wire [2:0] _0286_;
  wire [2:0] _0287_;
  wire [2:0] _0288_;
  wire [2:0] _0289_;
  wire [2:0] _0290_;
  wire [2:0] _0291_;
  wire [2:0] _0292_;
  wire [1:0] _0293_;
  wire [1:0] _0294_;
  wire _0295_;
  wire _0296_;
  wire _0297_;
  wire _0298_;
  wire _0299_;
  wire _0300_;
  wire _0301_;
  wire _0302_;
  wire _0303_;
  wire _0304_;
  wire _0305_;
  wire _0306_;
  wire _0307_;
  wire _0308_;
  wire _0309_;
  wire _0310_;
  wire _0311_;
  wire _0312_;
  wire _0313_;
  wire _0314_;
  wire _0315_;
  wire [31:0] _0316_;
  wire [31:0] _0317_;
  wire [31:0] _0318_;
  wire [31:0] _0319_;
  wire [31:0] _0320_;
  wire [31:0] _0321_;
  wire [31:0] _0322_;
  wire [31:0] _0323_;
  wire [31:0] _0324_;
  wire [31:0] _0325_;
  wire [31:0] _0326_;
  wire [31:0] _0327_;
  wire [31:0] _0328_;
  wire [31:0] _0329_;
  wire [31:0] _0330_;
  wire [31:0] _0331_;
  wire [31:0] _0332_;
  wire [31:0] _0333_;
  wire [31:0] _0334_;
  wire [31:0] _0335_;
  wire [31:0] _0336_;
  wire [31:0] _0337_;
  wire [31:0] _0338_;
  wire [31:0] _0339_;
  wire _0340_;
  wire _0341_;
  wire _0342_;
  wire _0343_;
  wire [31:0] _0344_;
  wire [31:0] _0345_;
  wire [31:0] _0346_;
  wire [31:0] _0347_;
  wire [31:0] _0348_;
  wire [31:0] _0349_;
  wire [31:0] _0350_;
  wire [31:0] _0351_;
  wire [31:0] _0352_;
  wire [31:0] _0353_;
  wire [31:0] _0354_;
  wire [31:0] _0355_;
  wire [31:0] _0356_;
  wire [31:0] _0357_;
  wire [31:0] _0358_;
  wire [31:0] _0359_;
  wire [31:0] _0360_;
  wire _0361_;
  wire _0362_;
  wire _0363_;
  wire _0364_;
  wire [31:0] _0365_;
  wire [31:0] _0366_;
  wire [31:0] _0367_;
  wire [31:0] _0368_;
  wire [31:0] _0369_;
  wire [31:0] _0370_;
  wire [31:0] _0371_;
  wire _0372_;
  wire _0373_;
  wire _0374_;
  wire _0375_;
  wire _0376_;
  wire _0377_;
  wire _0378_;
  wire [31:0] _0379_;
  wire [31:0] _0380_;
  wire [31:0] _0381_;
  wire [31:0] _0382_;
  wire [31:0] _0383_;
  wire [31:0] _0384_;
  wire [31:0] _0385_;
  wire [31:0] _0386_;
  wire [31:0] _0387_;
  wire [31:0] _0388_;
  wire [31:0] _0389_;
  wire [31:0] _0390_;
  wire [31:0] _0391_;
  wire [31:0] _0392_;
  wire [31:0] _0393_;
  wire [31:0] _0394_;
  wire _0395_;
  wire _0396_;
  wire [31:0] _0397_;
  wire [31:0] _0398_;
  wire [31:0] _0399_;
  wire [31:0] _0400_;
  wire [31:0] _0401_;
  wire [31:0] _0402_;
  wire _0403_;
  wire _0404_;
  wire _0405_;
  wire [31:0] _0406_;
  wire [31:0] _0407_;
  wire [31:0] _0408_;
  wire [31:0] _0409_;
  wire [31:0] _0410_;
  wire [31:0] _0411_;
  wire [31:0] _0412_;
  wire [31:0] _0413_;
  wire _0414_;
  wire [31:0] _0415_;
  wire [31:0] _0416_;
  wire [31:0] _0417_;
  wire [31:0] _0418_;
  wire [31:0] _0419_;
  wire [31:0] _0420_;
  wire [31:0] _0421_;
  wire _0422_;
  wire _0423_;
  wire [31:0] _0424_;
  wire [31:0] _0425_;
  wire [31:0] _0426_;
  wire _0427_;
  wire _0428_;
  wire [31:0] _0429_;
  wire [31:0] _0430_;
  wire [31:0] _0431_;
  wire [31:0] _0432_;
  wire [31:0] _0433_;
  wire [31:0] _0434_;
  wire [31:0] _0435_;
  wire [31:0] _0436_;
  wire _0437_;
  wire _0438_;
  wire _0439_;
  wire _0440_;
  wire _0441_;
  wire _0442_;
  wire _0443_;
  wire _0444_;
  wire _0445_;
  wire _0446_;
  wire _0447_;
  wire _0448_;
  wire _0449_;
  wire _0450_;
  wire _0451_;
  wire _0452_;
  wire _0453_;
  wire _0454_;
  wire _0455_;
  wire _0456_;
  wire _0457_;
  wire _0458_;
  wire _0459_;
  wire _0460_;
  wire _0461_;
  wire [31:0] _0462_;
  wire [31:0] _0463_;
  wire [31:0] _0464_;
  wire [31:0] _0465_;
  wire [31:0] _0466_;
  wire [31:0] _0467_;
  wire [31:0] _0468_;
  wire [31:0] _0469_;
  wire [31:0] _0470_;
  wire [31:0] _0471_;
  wire [31:0] _0472_;
  wire [31:0] _0473_;
  wire _0474_;
  wire _0475_;
  wire [31:0] _0476_;
  wire [31:0] _0477_;
  wire [31:0] _0478_;
  wire [31:0] _0479_;
  wire [31:0] _0480_;
  wire [31:0] _0481_;
  wire [31:0] _0482_;
  wire [31:0] _0483_;
  wire [31:0] _0484_;
  wire [31:0] _0485_;
  wire _0486_;
  wire _0487_;
  wire _0488_;
  wire [31:0] _0489_;
  wire [31:0] _0490_;
  wire [31:0] _0491_;
  wire [31:0] _0492_;
  wire _0493_;
  wire _0494_;
  wire _0495_;
  wire _0496_;
  wire [31:0] _0497_;
  wire [31:0] _0498_;
  wire [31:0] _0499_;
  wire [31:0] _0500_;
  wire _0501_;
  wire _0502_;
  wire _0503_;
  wire _0504_;
  wire _0505_;
  wire _0506_;
  wire _0507_;
  wire _0508_;
  wire _0509_;
  wire _0510_;
  wire _0511_;
  wire _0512_;
  wire _0513_;
  wire _0514_;
  wire _0515_;
  wire _0516_;
  wire [3:0] _0517_;
  wire [3:0] _0518_;
  wire _0519_;
  wire _0520_;
  wire _0521_;
  wire [3:0] _0522_;
  wire [3:0] _0523_;
  wire _0524_;
  wire _0525_;
  wire _0526_;
  wire _0527_;
  wire _0528_;
  wire _0529_;
  wire _0530_;
  wire _0531_;
  wire _0532_;
  wire _0533_;
  wire _0534_;
  wire _0535_;
  wire _0536_;
  wire _0537_;
  wire _0538_;
  wire _0539_;
  wire _0540_;
  wire _0541_;
  wire _0542_;
  wire _0543_;
  input clk_i;
  wire clk_i;
  output illegal_instr_o;
  wire illegal_instr_o;
  output illegal_instr_o_t0;
  wire illegal_instr_o_t0;
  input [31:0] instr_i;
  wire [31:0] instr_i;
  input [31:0] instr_i_t0;
  wire [31:0] instr_i_t0;
  output [31:0] instr_o;
  wire [31:0] instr_o;
  output [31:0] instr_o_t0;
  wire [31:0] instr_o_t0;
  output is_compressed_o;
  wire is_compressed_o;
  output is_compressed_o_t0;
  wire is_compressed_o_t0;
  input rst_ni;
  wire rst_ni;
  input valid_i;
  wire valid_i;
  input valid_i_t0;
  wire valid_i_t0;
  assign _0114_ = | { instr_i_t0[12], instr_i_t0[6:5] };
  assign _0115_ = | instr_i_t0[11:10];
  assign _0111_ = | instr_i_t0[1:0];
  assign _0083_ = ~ instr_i_t0[11:7];
  assign _0094_ = ~ { instr_i_t0[12], instr_i_t0[6:5] };
  assign _0095_ = ~ instr_i_t0[11:10];
  assign _0100_ = ~ instr_i_t0[15:13];
  assign _0086_ = ~ instr_i_t0[1:0];
  assign _0244_ = instr_i[11:7] & _0083_;
  assign _0268_ = { instr_i[12], instr_i[6:5] } & _0094_;
  assign _0276_ = instr_i[11:10] & _0095_;
  assign _0285_ = instr_i[15:13] & _0100_;
  assign _0248_ = instr_i[1:0] & _0086_;
  assign _0245_ = 5'h02 & _0083_;
  assign _0269_ = 3'h4 & _0094_;
  assign _0270_ = 3'h5 & _0094_;
  assign _0271_ = 3'h6 & _0094_;
  assign _0272_ = 3'h7 & _0094_;
  assign _0273_ = 3'h3 & _0094_;
  assign _0274_ = 3'h2 & _0094_;
  assign _0275_ = 3'h1 & _0094_;
  assign _0277_ = 2'h3 & _0095_;
  assign _0278_ = 2'h2 & _0095_;
  assign _0286_ = 3'h1 & _0100_;
  assign _0287_ = 3'h3 & _0100_;
  assign _0288_ = 3'h4 & _0100_;
  assign _0289_ = 3'h5 & _0100_;
  assign _0290_ = 3'h7 & _0100_;
  assign _0291_ = 3'h6 & _0100_;
  assign _0292_ = 3'h2 & _0100_;
  assign _0293_ = 2'h1 & _0086_;
  assign _0249_ = 2'h3 & _0086_;
  assign _0294_ = 2'h2 & _0086_;
  assign _0437_ = _0244_ == _0245_;
  assign _0439_ = _0268_ == _0269_;
  assign _0440_ = _0268_ == _0270_;
  assign _0441_ = _0268_ == _0271_;
  assign _0442_ = _0268_ == _0272_;
  assign _0443_ = _0268_ == _0273_;
  assign _0444_ = _0268_ == _0274_;
  assign _0445_ = _0268_ == _0275_;
  assign _0446_ = _0276_ == _0277_;
  assign _0447_ = _0276_ == _0278_;
  assign _0448_ = _0285_ == _0286_;
  assign _0449_ = _0285_ == _0287_;
  assign _0450_ = _0285_ == _0288_;
  assign _0451_ = _0285_ == _0289_;
  assign _0452_ = _0285_ == _0290_;
  assign _0453_ = _0285_ == _0291_;
  assign _0454_ = _0285_ == _0292_;
  assign _0455_ = _0248_ == _0293_;
  assign _0438_ = _0248_ == _0249_;
  assign _0456_ = _0248_ == _0294_;
  assign _0503_ = _0437_ & _0108_;
  assign is_compressed_o_t0 = _0438_ & _0111_;
  assign _0523_[0] = _0439_ & _0114_;
  assign _0523_[1] = _0440_ & _0114_;
  assign _0523_[2] = _0441_ & _0114_;
  assign _0523_[3] = _0442_ & _0114_;
  assign _0526_ = _0443_ & _0114_;
  assign _0528_ = _0444_ & _0114_;
  assign _0530_ = _0445_ & _0114_;
  assign _0532_ = _0446_ & _0115_;
  assign _0536_ = _0447_ & _0115_;
  assign _0518_[0] = _0448_ & _0119_;
  assign _0518_[1] = _0449_ & _0119_;
  assign _0510_ = _0450_ & _0119_;
  assign _0518_[2] = _0451_ & _0119_;
  assign _0518_[3] = _0452_ & _0119_;
  assign _0521_ = _0453_ & _0119_;
  assign _0514_ = _0454_ & _0119_;
  assign _0534_ = _0455_ & _0111_;
  assign _0512_ = _0456_ & _0111_;
  assign _0104_ = | { _0514_, _0521_ };
  assign _0105_ = | { _0514_, _0521_, _0516_, _0518_[3:2], _0518_[0] };
  assign _0106_ = | { _0521_, _0518_[3], _0518_[1], _0510_ };
  assign _0107_ = | instr_i_t0[12:5];
  assign _0109_ = | { instr_i_t0[12], instr_i_t0[6:2] };
  assign _0108_ = | instr_i_t0[11:7];
  assign _0110_ = | instr_i_t0[6:2];
  assign _0112_ = | _0518_;
  assign _0113_ = | _0523_;
  assign _0116_ = | { _0521_, _0518_[3] };
  assign _0117_ = | { _0518_[2], _0518_[0] };
  assign _0118_ = | { _0518_, _0510_ };
  assign _0119_ = | instr_i_t0[15:13];
  assign _0045_ = ~ { _0521_, _0514_ };
  assign _0046_ = ~ { _0521_, _0518_[3:2], _0518_[0], _0516_, _0514_ };
  assign _0054_ = ~ { _0521_, _0518_[3], _0518_[1], _0510_ };
  assign _0082_ = ~ instr_i_t0[12:5];
  assign _0084_ = ~ { instr_i_t0[12], instr_i_t0[6:2] };
  assign _0085_ = ~ instr_i_t0[6:2];
  assign _0092_ = ~ _0518_;
  assign _0093_ = ~ _0523_;
  assign _0097_ = ~ { _0521_, _0518_[3] };
  assign _0098_ = ~ { _0518_[2], _0518_[0] };
  assign _0099_ = ~ { _0518_, _0510_ };
  assign _0133_ = { _0520_, _0513_ } & _0045_;
  assign _0134_ = { _0520_, _0517_[3:2], _0517_[0], _0515_, _0513_ } & _0046_;
  assign _0147_ = { _0520_, _0517_[3], _0517_[1], _0509_ } & _0054_;
  assign _0243_ = instr_i[12:5] & _0082_;
  assign _0246_ = { instr_i[12], instr_i[6:2] } & _0084_;
  assign _0247_ = instr_i[6:2] & _0085_;
  assign _0266_ = _0517_ & _0092_;
  assign _0267_ = _0522_ & _0093_;
  assign _0282_ = { _0520_, _0517_[3] } & _0097_;
  assign _0283_ = { _0517_[2], _0517_[0] } & _0098_;
  assign _0284_ = { _0517_, _0509_ } & _0099_;
  assign _0120_ = ! _0133_;
  assign _0121_ = ! _0134_;
  assign _0122_ = ! _0147_;
  assign _0123_ = ! _0243_;
  assign _0124_ = ! _0246_;
  assign _0125_ = ! _0244_;
  assign _0126_ = ! _0247_;
  assign _0127_ = ! _0266_;
  assign _0128_ = ! _0267_;
  assign _0129_ = ! _0282_;
  assign _0130_ = ! _0283_;
  assign _0131_ = ! _0284_;
  assign _0132_ = ! _0285_;
  assign _0042_ = _0120_ & _0104_;
  assign _0044_ = _0121_ & _0105_;
  assign _0103_ = _0122_ & _0106_;
  assign _0016_ = _0123_ & _0107_;
  assign _0024_ = _0124_ & _0109_;
  assign _0004_ = _0125_ & _0108_;
  assign _0507_ = _0126_ & _0110_;
  assign _0148_ = _0127_ & _0112_;
  assign _0034_ = _0128_ & _0113_;
  assign _0538_ = _0129_ & _0116_;
  assign _0540_ = _0130_ & _0117_;
  assign _0542_ = _0131_ & _0118_;
  assign _0516_ = _0132_ & _0119_;
  assign _0048_ = ~ _0519_;
  assign _0055_ = ~ _0513_;
  assign _0057_ = ~ _0295_;
  assign _0058_ = ~ { _0519_, _0519_, _0519_, _0519_, _0519_, _0519_, _0519_, _0519_, _0519_, _0519_, _0519_, _0519_, _0519_, _0519_, _0519_, _0519_, _0519_, _0519_, _0519_, _0519_, _0519_, _0519_, _0519_, _0519_, _0519_, _0519_, _0519_, _0519_, _0519_, _0519_, _0519_, _0519_ };
  assign _0061_ = ~ { _0295_, _0295_, _0295_, _0295_, _0295_, _0295_, _0295_, _0295_, _0295_, _0295_, _0295_, _0295_, _0295_, _0295_, _0295_, _0295_, _0295_, _0295_, _0295_, _0295_, _0295_, _0295_, _0295_, _0295_, _0295_, _0295_, _0295_, _0295_, _0295_, _0295_, _0295_, _0295_ };
  assign _0062_ = ~ { _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_ };
  assign _0063_ = ~ { _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_ };
  assign _0064_ = ~ { _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_ };
  assign _0065_ = ~ { _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_ };
  assign _0050_ = ~ _0524_;
  assign _0066_ = ~ _0535_;
  assign _0067_ = ~ _0531_;
  assign _0068_ = ~ { _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_ };
  assign _0069_ = ~ { _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_ };
  assign _0060_ = ~ { _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_ };
  assign _0070_ = ~ { _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_ };
  assign _0071_ = ~ { _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_ };
  assign _0072_ = ~ { _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_ };
  assign _0056_ = ~ _0509_;
  assign _0073_ = ~ _0043_;
  assign _0074_ = ~ _0041_;
  assign _0051_ = ~ _0541_;
  assign _0075_ = ~ { _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_ };
  assign _0059_ = ~ { _0513_, _0513_, _0513_, _0513_, _0513_, _0513_, _0513_, _0513_, _0513_, _0513_, _0513_, _0513_, _0513_, _0513_, _0513_, _0513_, _0513_, _0513_, _0513_, _0513_, _0513_, _0513_, _0513_, _0513_, _0513_, _0513_, _0513_, _0513_, _0513_, _0513_, _0513_, _0513_ };
  assign _0076_ = ~ { _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_ };
  assign _0053_ = ~ _0543_;
  assign _0077_ = ~ _0533_;
  assign _0078_ = ~ _0301_;
  assign _0079_ = ~ { _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_ };
  assign _0080_ = ~ { _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_ };
  assign _0081_ = ~ { _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_ };
  assign _0087_ = ~ { _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_ };
  assign _0088_ = ~ { _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_ };
  assign _0089_ = ~ _0506_;
  assign _0091_ = ~ { instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12] };
  assign _0090_ = ~ instr_i[12];
  assign _0096_ = ~ { _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_ };
  assign _0307_ = _0514_ | _0055_;
  assign _0313_ = _0296_ | _0057_;
  assign _0316_ = { _0148_, _0148_, _0148_, _0148_, _0148_, _0148_, _0148_, _0148_, _0148_, _0148_, _0148_, _0148_, _0148_, _0148_, _0148_, _0148_, _0148_, _0148_, _0148_, _0148_, _0148_, _0148_, _0148_, _0148_, _0148_, _0148_, _0148_, _0148_, _0148_, _0148_, _0148_, _0148_ } | _0058_;
  assign _0325_ = { _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_ } | _0061_;
  assign _0328_ = { _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_ } | _0062_;
  assign _0331_ = { _0530_, _0530_, _0530_, _0530_, _0530_, _0530_, _0530_, _0530_, _0530_, _0530_, _0530_, _0530_, _0530_, _0530_, _0530_, _0530_, _0530_, _0530_, _0530_, _0530_, _0530_, _0530_, _0530_, _0530_, _0530_, _0530_, _0530_, _0530_, _0530_, _0530_, _0530_, _0530_ } | _0063_;
  assign _0334_ = { _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_ } | _0064_;
  assign _0337_ = { _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_ } | _0065_;
  assign _0340_ = _0536_ | _0066_;
  assign _0341_ = _0532_ | _0067_;
  assign _0344_ = { _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_ } | _0068_;
  assign _0347_ = { _0532_, _0532_, _0532_, _0532_, _0532_, _0532_, _0532_, _0532_, _0532_, _0532_, _0532_, _0532_, _0532_, _0532_, _0532_, _0532_, _0532_, _0532_, _0532_, _0532_, _0532_, _0532_, _0532_, _0532_, _0532_, _0532_, _0532_, _0532_, _0532_, _0532_, _0532_, _0532_ } | _0069_;
  assign _0322_ = { _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_ } | _0060_;
  assign _0351_ = { _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_ } | _0070_;
  assign _0354_ = { _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_ } | _0071_;
  assign _0358_ = { _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_ } | _0072_;
  assign _0310_ = _0510_ | _0056_;
  assign _0362_ = _0044_ | _0073_;
  assign _0363_ = _0042_ | _0074_;
  assign _0364_ = _0542_ | _0051_;
  assign _0365_ = { _0542_, _0542_, _0542_, _0542_, _0542_, _0542_, _0542_, _0542_, _0542_, _0542_, _0542_, _0542_, _0542_, _0542_, _0542_, _0542_, _0542_, _0542_, _0542_, _0542_, _0542_, _0542_, _0542_, _0542_, _0542_, _0542_, _0542_, _0542_, _0542_, _0542_, _0542_, _0542_ } | _0075_;
  assign _0319_ = { _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_ } | _0059_;
  assign _0369_ = { _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_ } | _0076_;
  assign _0372_ = is_compressed_o_t0 | _0053_;
  assign _0373_ = _0534_ | _0077_;
  assign _0376_ = _0302_ | _0078_;
  assign _0379_ = { is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0 } | _0079_;
  assign _0382_ = { _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_ } | _0080_;
  assign _0385_ = { _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_ } | _0081_;
  assign _0388_ = { _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_ } | _0087_;
  assign _0391_ = { _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_ } | _0088_;
  assign _0395_ = _0507_ | _0089_;
  assign _0397_ = { instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12] } | _0091_;
  assign _0396_ = instr_i_t0[12] | _0090_;
  assign _0400_ = { _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_ } | _0096_;
  assign _0308_ = _0514_ | _0513_;
  assign _0314_ = _0296_ | _0295_;
  assign _0317_ = { _0148_, _0148_, _0148_, _0148_, _0148_, _0148_, _0148_, _0148_, _0148_, _0148_, _0148_, _0148_, _0148_, _0148_, _0148_, _0148_, _0148_, _0148_, _0148_, _0148_, _0148_, _0148_, _0148_, _0148_, _0148_, _0148_, _0148_, _0148_, _0148_, _0148_, _0148_, _0148_ } | { _0519_, _0519_, _0519_, _0519_, _0519_, _0519_, _0519_, _0519_, _0519_, _0519_, _0519_, _0519_, _0519_, _0519_, _0519_, _0519_, _0519_, _0519_, _0519_, _0519_, _0519_, _0519_, _0519_, _0519_, _0519_, _0519_, _0519_, _0519_, _0519_, _0519_, _0519_, _0519_ };
  assign _0326_ = { _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_ } | { _0295_, _0295_, _0295_, _0295_, _0295_, _0295_, _0295_, _0295_, _0295_, _0295_, _0295_, _0295_, _0295_, _0295_, _0295_, _0295_, _0295_, _0295_, _0295_, _0295_, _0295_, _0295_, _0295_, _0295_, _0295_, _0295_, _0295_, _0295_, _0295_, _0295_, _0295_, _0295_ };
  assign _0329_ = { _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_ } | { _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_ };
  assign _0332_ = { _0530_, _0530_, _0530_, _0530_, _0530_, _0530_, _0530_, _0530_, _0530_, _0530_, _0530_, _0530_, _0530_, _0530_, _0530_, _0530_, _0530_, _0530_, _0530_, _0530_, _0530_, _0530_, _0530_, _0530_, _0530_, _0530_, _0530_, _0530_, _0530_, _0530_, _0530_, _0530_ } | { _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_ };
  assign _0335_ = { _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_ } | { _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_ };
  assign _0338_ = { _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_ } | { _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_ };
  assign _0342_ = _0532_ | _0531_;
  assign _0345_ = { _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_ } | { _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_ };
  assign _0348_ = { _0532_, _0532_, _0532_, _0532_, _0532_, _0532_, _0532_, _0532_, _0532_, _0532_, _0532_, _0532_, _0532_, _0532_, _0532_, _0532_, _0532_, _0532_, _0532_, _0532_, _0532_, _0532_, _0532_, _0532_, _0532_, _0532_, _0532_, _0532_, _0532_, _0532_, _0532_, _0532_ } | { _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_ };
  assign _0323_ = { _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_ } | { _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_ };
  assign _0352_ = { _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_ } | { _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_ };
  assign _0355_ = { _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_ } | { _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_ };
  assign _0359_ = { _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_ } | { _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_ };
  assign _0311_ = _0510_ | _0509_;
  assign _0366_ = { _0542_, _0542_, _0542_, _0542_, _0542_, _0542_, _0542_, _0542_, _0542_, _0542_, _0542_, _0542_, _0542_, _0542_, _0542_, _0542_, _0542_, _0542_, _0542_, _0542_, _0542_, _0542_, _0542_, _0542_, _0542_, _0542_, _0542_, _0542_, _0542_, _0542_, _0542_, _0542_ } | { _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_ };
  assign _0320_ = { _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_ } | { _0513_, _0513_, _0513_, _0513_, _0513_, _0513_, _0513_, _0513_, _0513_, _0513_, _0513_, _0513_, _0513_, _0513_, _0513_, _0513_, _0513_, _0513_, _0513_, _0513_, _0513_, _0513_, _0513_, _0513_, _0513_, _0513_, _0513_, _0513_, _0513_, _0513_, _0513_, _0513_ };
  assign _0370_ = { _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_ } | { _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_ };
  assign _0374_ = _0534_ | _0533_;
  assign _0377_ = _0302_ | _0301_;
  assign _0380_ = { is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0 } | { _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_ };
  assign _0383_ = { _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_ } | { _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_ };
  assign _0386_ = { _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_ } | { _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_ };
  assign _0389_ = { _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_ } | { _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_ };
  assign _0392_ = { _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_ } | { _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_ };
  assign _0398_ = { instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12] } | { instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12] };
  assign _0401_ = { _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_ } | { _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_ };
  assign _0149_ = instr_i_t0[12] & _0307_;
  assign _0152_ = _0459_ & _0310_;
  assign _0155_ = _0461_ & _0313_;
  assign _0158_ = { 4'h0, instr_i_t0[8:7], instr_i_t0[12], instr_i_t0[6:2], 8'h00, instr_i_t0[11:9], 9'h000 } & _0316_;
  assign _0161_ = { 7'h00, instr_i_t0[6:2], instr_i_t0[11:7], 3'h0, instr_i_t0[11:7], 7'h00 } & _0319_;
  assign _0164_ = _0465_ & _0322_;
  assign _0167_ = _0467_ & _0325_;
  assign _0170_ = { 9'h000, instr_i_t0[4:2], 2'h0, instr_i_t0[9:7], 5'h00, instr_i_t0[9:7], 7'h00 } & _0328_;
  assign _0173_ = { 9'h000, instr_i_t0[4:2], 2'h0, instr_i_t0[9:7], 5'h00, instr_i_t0[9:7], 7'h00 } & _0331_;
  assign _0176_ = _0471_ & _0334_;
  assign _0179_ = _0473_ & _0337_;
  assign _0182_ = instr_i_t0[12] & _0340_;
  assign _0184_ = _0475_ & _0341_;
  assign _0187_ = { 1'h0, instr_i_t0[10], 5'h00, instr_i_t0[6:2], 2'h0, instr_i_t0[9:7], 5'h00, instr_i_t0[9:7], 7'h00 } & _0344_;
  assign _0190_ = _0477_ & _0347_;
  assign _0193_ = _0022_ & _0322_;
  assign _0196_ = _0479_ & _0351_;
  assign _0199_ = { instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[6:2], instr_i_t0[11:7], 3'h0, instr_i_t0[11:7], 7'h00 } & _0354_;
  assign _0202_ = _0483_ & _0319_;
  assign _0205_ = _0485_ & _0358_;
  assign _0208_ = _0024_ & _0310_;
  assign _0211_ = _0486_ & _0362_;
  assign _0213_ = _0016_ & _0363_;
  assign _0215_ = _0488_ & _0364_;
  assign _0217_ = { 5'h00, instr_i_t0[5], instr_i_t0[12], 2'h0, instr_i_t0[4:2], 2'h0, instr_i_t0[9:7], 3'h0, instr_i_t0[11:10], instr_i_t0[6], 9'h000 } & _0365_;
  assign _0220_ = { 2'h0, instr_i_t0[10:7], instr_i_t0[12:11], instr_i_t0[5], instr_i_t0[6], 12'h000, instr_i_t0[4:2], 7'h00 } & _0319_;
  assign _0223_ = _0492_ & _0369_;
  assign _0226_ = _0038_ & _0372_;
  assign _0228_ = _0012_ & _0373_;
  assign _0231_ = _0496_ & _0376_;
  assign _0234_ = _0032_ & _0379_;
  assign _0237_ = _0014_ & _0382_;
  assign _0240_ = _0500_ & _0385_;
  assign _0250_ = { 12'h000, instr_i_t0[11:7], 15'h0000 } & _0388_;
  assign _0253_ = _0006_ & _0391_;
  assign _0256_ = { 12'h000, instr_i_t0[11:7], 15'h0000 } & _0391_;
  assign _0259_ = _0004_ & _0395_;
  assign _0261_ = _0010_ & _0396_;
  assign _0263_ = _0040_ & _0397_;
  assign _0279_ = { instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[6:2], instr_i_t0[11:7], 7'h00 } & _0400_;
  assign _0150_ = _0004_ & _0308_;
  assign _0153_ = _0008_ & _0311_;
  assign _0156_ = _0148_ & _0314_;
  assign _0159_ = instr_i_t0 & _0317_;
  assign _0162_ = { 4'h0, instr_i_t0[3:2], instr_i_t0[12], instr_i_t0[6:4], 10'h000, instr_i_t0[11:7], 7'h00 } & _0320_;
  assign _0165_ = _0036_ & _0323_;
  assign _0168_ = _0463_ & _0326_;
  assign _0171_ = instr_i_t0 & _0329_;
  assign _0174_ = { 9'h000, instr_i_t0[4:2], 2'h0, instr_i_t0[9:7], 5'h00, instr_i_t0[9:7], 7'h00 } & _0332_;
  assign _0177_ = { 9'h000, instr_i_t0[4:2], 2'h0, instr_i_t0[9:7], 5'h00, instr_i_t0[9:7], 7'h00 } & _0335_;
  assign _0180_ = _0469_ & _0338_;
  assign _0185_ = _0034_ & _0342_;
  assign _0188_ = { instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[6:2], 2'h0, instr_i_t0[9:7], 5'h00, instr_i_t0[9:7], 7'h00 } & _0345_;
  assign _0191_ = _0030_ & _0348_;
  assign _0194_ = _0026_ & _0323_;
  assign _0197_ = { instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[6:5], instr_i_t0[2], 7'h00, instr_i_t0[9:7], 2'h0, instr_i_t0[13], instr_i_t0[11:10], instr_i_t0[4:3], instr_i_t0[12], 7'h00 } & _0352_;
  assign _0200_ = { instr_i_t0[12], instr_i_t0[8], instr_i_t0[10:9], instr_i_t0[6], instr_i_t0[7], instr_i_t0[2], instr_i_t0[11], instr_i_t0[5:3], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], 4'h0, instr_i_t0[15], 7'h00 } & _0355_;
  assign _0203_ = { instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[6:2], 8'h00, instr_i_t0[11:7], 7'h00 } & _0320_;
  assign _0206_ = _0481_ & _0359_;
  assign _0209_ = _0028_ & _0311_;
  assign _0218_ = instr_i_t0 & _0366_;
  assign _0221_ = { 5'h00, instr_i_t0[5], instr_i_t0[12:10], instr_i_t0[6], 4'h0, instr_i_t0[9:7], 5'h00, instr_i_t0[4:2], 7'h00 } & _0320_;
  assign _0224_ = _0490_ & _0370_;
  assign _0229_ = _0020_ & _0374_;
  assign _0232_ = _0494_ & _0377_;
  assign _0235_ = instr_i_t0 & _0380_;
  assign _0238_ = _0018_ & _0383_;
  assign _0241_ = _0498_ & _0386_;
  assign _0251_ = 32'd0 & _0389_;
  assign _0254_ = { 7'h00, instr_i_t0[6:2], instr_i_t0[11:7], 3'h0, instr_i_t0[11:7], 7'h00 } & _0392_;
  assign _0257_ = { 7'h00, instr_i_t0[6:2], 8'h00, instr_i_t0[11:7], 7'h00 } & _0392_;
  assign _0264_ = _0002_ & _0398_;
  assign _0280_ = { instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[4:3], instr_i_t0[5], instr_i_t0[2], instr_i_t0[6], 24'h000000 } & _0401_;
  assign _0309_ = _0149_ | _0150_;
  assign _0312_ = _0152_ | _0153_;
  assign _0315_ = _0155_ | _0156_;
  assign _0318_ = _0158_ | _0159_;
  assign _0321_ = _0161_ | _0162_;
  assign _0324_ = _0164_ | _0165_;
  assign _0327_ = _0167_ | _0168_;
  assign _0330_ = _0170_ | _0171_;
  assign _0333_ = _0173_ | _0174_;
  assign _0336_ = _0176_ | _0177_;
  assign _0339_ = _0179_ | _0180_;
  assign _0343_ = _0184_ | _0185_;
  assign _0346_ = _0187_ | _0188_;
  assign _0349_ = _0190_ | _0191_;
  assign _0350_ = _0193_ | _0194_;
  assign _0353_ = _0196_ | _0197_;
  assign _0356_ = _0199_ | _0200_;
  assign _0357_ = _0202_ | _0203_;
  assign _0360_ = _0205_ | _0206_;
  assign _0361_ = _0208_ | _0209_;
  assign _0367_ = _0217_ | _0218_;
  assign _0368_ = _0220_ | _0221_;
  assign _0371_ = _0223_ | _0224_;
  assign _0375_ = _0228_ | _0229_;
  assign _0378_ = _0231_ | _0232_;
  assign _0381_ = _0234_ | _0235_;
  assign _0384_ = _0237_ | _0238_;
  assign _0387_ = _0240_ | _0241_;
  assign _0390_ = _0250_ | _0251_;
  assign _0393_ = _0253_ | _0254_;
  assign _0394_ = _0256_ | _0257_;
  assign _0399_ = _0263_ | _0264_;
  assign _0402_ = _0279_ | _0280_;
  assign _0403_ = _0000_ ^ _0003_;
  assign _0404_ = _0458_ ^ _0007_;
  assign _0405_ = _0460_ ^ _0457_;
  assign _0406_ = { 4'h0, instr_i[8:7], instr_i[12], instr_i[6:2], 8'h12, instr_i[11:9], 9'h023 } ^ instr_i;
  assign _0407_ = { 7'h00, instr_i[6:2], instr_i[11:7], 3'h1, instr_i[11:7], 7'h13 } ^ { 4'h0, instr_i[3:2], instr_i[12], instr_i[6:4], 10'h012, instr_i[11:7], 7'h03 };
  assign _0408_ = _0464_ ^ _0035_;
  assign _0409_ = _0466_ ^ _0462_;
  assign _0410_ = { 9'h001, instr_i[4:2], 2'h1, instr_i[9:7], 5'h1d, instr_i[9:7], 7'h33 } ^ instr_i;
  assign _0411_ = { 9'h081, instr_i[4:2], 2'h1, instr_i[9:7], 5'h01, instr_i[9:7], 7'h33 } ^ { 9'h001, instr_i[4:2], 2'h1, instr_i[9:7], 5'h11, instr_i[9:7], 7'h33 };
  assign _0412_ = _0470_ ^ { 9'h001, instr_i[4:2], 2'h1, instr_i[9:7], 5'h19, instr_i[9:7], 7'h33 };
  assign _0413_ = _0472_ ^ _0468_;
  assign _0414_ = _0474_ ^ _0033_;
  assign _0415_ = { 1'h0, instr_i[10], 5'h00, instr_i[6:2], 2'h1, instr_i[9:7], 5'h15, instr_i[9:7], 7'h13 } ^ { instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[6:2], 2'h1, instr_i[9:7], 5'h1d, instr_i[9:7], 7'h13 };
  assign _0416_ = _0476_ ^ _0029_;
  assign _0417_ = _0021_ ^ _0025_;
  assign _0418_ = _0478_ ^ { instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[6:5], instr_i[2], 7'h01, instr_i[9:7], 2'h0, instr_i[13], instr_i[11:10], instr_i[4:3], instr_i[12], 7'h63 };
  assign _0419_ = { instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[6:2], instr_i[11:7], 3'h0, instr_i[11:7], 7'h13 } ^ { instr_i[12], instr_i[8], instr_i[10:9], instr_i[6], instr_i[7], instr_i[2], instr_i[11], instr_i[5:3], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], 4'h0, _0508_, 7'h6f };
  assign _0420_ = _0482_ ^ { instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[6:2], 8'h00, instr_i[11:7], 7'h13 };
  assign _0421_ = _0484_ ^ _0480_;
  assign _0422_ = _0023_ ^ _0027_;
  assign _0424_ = { 5'h00, instr_i[5], instr_i[12], 2'h1, instr_i[4:2], 2'h1, instr_i[9:7], 3'h2, instr_i[11:10], instr_i[6], 9'h023 } ^ instr_i;
  assign _0425_ = { 2'h0, instr_i[10:7], instr_i[12:11], instr_i[5], instr_i[6], 12'h041, instr_i[4:2], 7'h13 } ^ { 5'h00, instr_i[5], instr_i[12:10], instr_i[6], 4'h1, instr_i[9:7], 5'h09, instr_i[4:2], 7'h03 };
  assign _0426_ = _0491_ ^ _0489_;
  assign _0427_ = _0011_ ^ _0019_;
  assign _0428_ = _0495_ ^ _0493_;
  assign _0429_ = _0031_ ^ instr_i;
  assign _0430_ = _0013_ ^ _0017_;
  assign _0431_ = _0499_ ^ _0497_;
  assign _0432_ = { 12'h000, instr_i[11:7], 15'h00e7 } ^ 32'd1048691;
  assign _0433_ = _0005_ ^ { 7'h00, instr_i[6:2], instr_i[11:7], 3'h0, instr_i[11:7], 7'h33 };
  assign _0434_ = { 12'h000, instr_i[11:7], 15'h0067 } ^ { 7'h00, instr_i[6:2], 8'h00, instr_i[11:7], 7'h33 };
  assign _0435_ = _0039_ ^ _0001_;
  assign _0436_ = { instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[6:2], instr_i[11:7], 7'h37 } ^ { instr_i[12], instr_i[12], instr_i[12], instr_i[4:3], instr_i[5], instr_i[2], instr_i[6], 24'h010113 };
  assign _0151_ = _0514_ & _0403_;
  assign _0154_ = _0510_ & _0404_;
  assign _0157_ = _0296_ & _0405_;
  assign _0160_ = { _0148_, _0148_, _0148_, _0148_, _0148_, _0148_, _0148_, _0148_, _0148_, _0148_, _0148_, _0148_, _0148_, _0148_, _0148_, _0148_, _0148_, _0148_, _0148_, _0148_, _0148_, _0148_, _0148_, _0148_, _0148_, _0148_, _0148_, _0148_, _0148_, _0148_, _0148_, _0148_ } & _0406_;
  assign _0163_ = { _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_ } & _0407_;
  assign _0166_ = { _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_ } & _0408_;
  assign _0169_ = { _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_ } & _0409_;
  assign _0172_ = { _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_ } & _0410_;
  assign _0175_ = { _0530_, _0530_, _0530_, _0530_, _0530_, _0530_, _0530_, _0530_, _0530_, _0530_, _0530_, _0530_, _0530_, _0530_, _0530_, _0530_, _0530_, _0530_, _0530_, _0530_, _0530_, _0530_, _0530_, _0530_, _0530_, _0530_, _0530_, _0530_, _0530_, _0530_, _0530_, _0530_ } & _0411_;
  assign _0178_ = { _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_ } & _0412_;
  assign _0181_ = { _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_ } & _0413_;
  assign _0183_ = _0536_ & _0000_;
  assign _0186_ = _0532_ & _0414_;
  assign _0189_ = { _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_ } & _0415_;
  assign _0192_ = { _0532_, _0532_, _0532_, _0532_, _0532_, _0532_, _0532_, _0532_, _0532_, _0532_, _0532_, _0532_, _0532_, _0532_, _0532_, _0532_, _0532_, _0532_, _0532_, _0532_, _0532_, _0532_, _0532_, _0532_, _0532_, _0532_, _0532_, _0532_, _0532_, _0532_, _0532_, _0532_ } & _0416_;
  assign _0195_ = { _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_ } & _0417_;
  assign _0198_ = { _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_ } & _0418_;
  assign _0201_ = { _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_, _0540_ } & _0419_;
  assign _0204_ = { _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_ } & _0420_;
  assign _0207_ = { _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_ } & _0421_;
  assign _0210_ = _0510_ & _0422_;
  assign _0212_ = _0044_ & _0423_;
  assign _0214_ = _0042_ & _0015_;
  assign _0216_ = _0542_ & _0101_;
  assign _0219_ = { _0542_, _0542_, _0542_, _0542_, _0542_, _0542_, _0542_, _0542_, _0542_, _0542_, _0542_, _0542_, _0542_, _0542_, _0542_, _0542_, _0542_, _0542_, _0542_, _0542_, _0542_, _0542_, _0542_, _0542_, _0542_, _0542_, _0542_, _0542_, _0542_, _0542_, _0542_, _0542_ } & _0424_;
  assign _0222_ = { _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_ } & _0425_;
  assign _0225_ = { _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_ } & _0426_;
  assign _0227_ = is_compressed_o_t0 & _0037_;
  assign _0230_ = _0534_ & _0427_;
  assign _0233_ = _0302_ & _0428_;
  assign _0236_ = { is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0 } & _0429_;
  assign _0239_ = { _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_ } & _0430_;
  assign _0242_ = { _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_ } & _0431_;
  assign _0252_ = { _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_ } & _0432_;
  assign _0255_ = { _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_ } & _0433_;
  assign _0258_ = { _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_ } & _0434_;
  assign _0260_ = _0507_ & _0003_;
  assign _0262_ = instr_i_t0[12] & _0009_;
  assign _0265_ = { instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12] } & _0435_;
  assign _0281_ = { _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_ } & _0436_;
  assign _0459_ = _0151_ | _0309_;
  assign _0461_ = _0154_ | _0312_;
  assign _0038_ = _0157_ | _0315_;
  assign _0463_ = _0160_ | _0318_;
  assign _0465_ = _0163_ | _0321_;
  assign _0467_ = _0166_ | _0324_;
  assign _0032_ = _0169_ | _0327_;
  assign _0469_ = _0172_ | _0330_;
  assign _0471_ = _0175_ | _0333_;
  assign _0473_ = _0178_ | _0336_;
  assign _0030_ = _0181_ | _0339_;
  assign _0475_ = _0183_ | _0182_;
  assign _0028_ = _0186_ | _0343_;
  assign _0477_ = _0189_ | _0346_;
  assign _0026_ = _0192_ | _0349_;
  assign _0479_ = _0195_ | _0350_;
  assign _0481_ = _0198_ | _0353_;
  assign _0483_ = _0201_ | _0356_;
  assign _0485_ = _0204_ | _0357_;
  assign _0018_ = _0207_ | _0360_;
  assign _0486_ = _0210_ | _0361_;
  assign _0020_ = _0212_ | _0211_;
  assign _0488_ = _0214_ | _0213_;
  assign _0012_ = _0216_ | _0215_;
  assign _0490_ = _0219_ | _0367_;
  assign _0492_ = _0222_ | _0368_;
  assign _0014_ = _0225_ | _0371_;
  assign _0494_ = _0227_ | _0226_;
  assign _0496_ = _0230_ | _0375_;
  assign illegal_instr_o_t0 = _0233_ | _0378_;
  assign _0498_ = _0236_ | _0381_;
  assign _0500_ = _0239_ | _0384_;
  assign instr_o_t0 = _0242_ | _0387_;
  assign _0006_ = _0252_ | _0390_;
  assign _0002_ = _0255_ | _0393_;
  assign _0040_ = _0258_ | _0394_;
  assign _0010_ = _0260_ | _0259_;
  assign _0008_ = _0262_ | _0261_;
  assign _0036_ = _0265_ | _0399_;
  assign _0022_ = _0281_ | _0402_;
  assign _0101_ = ~ _0487_;
  assign _0041_ = | { _0520_, _0513_ };
  assign _0043_ = | { _0520_, _0517_[3:2], _0517_[0], _0515_, _0513_ };
  assign _0049_ = ~ _0525_;
  assign _0047_ = ~ _0520_;
  assign _0052_ = ~ _0511_;
  assign _0135_ = _0521_ & _0048_;
  assign _0138_ = _0526_ & _0050_;
  assign _0141_ = _0521_ & _0051_;
  assign _0144_ = _0512_ & _0053_;
  assign _0136_ = _0148_ & _0047_;
  assign _0139_ = _0034_ & _0049_;
  assign _0142_ = _0542_ & _0047_;
  assign _0145_ = is_compressed_o_t0 & _0052_;
  assign _0137_ = _0521_ & _0148_;
  assign _0140_ = _0526_ & _0034_;
  assign _0143_ = _0521_ & _0542_;
  assign _0146_ = _0512_ & is_compressed_o_t0;
  assign _0303_ = _0135_ | _0136_;
  assign _0304_ = _0138_ | _0139_;
  assign _0305_ = _0141_ | _0142_;
  assign _0306_ = _0144_ | _0145_;
  assign _0296_ = _0303_ | _0137_;
  assign _0298_ = _0304_ | _0140_;
  assign _0300_ = _0305_ | _0143_;
  assign _0302_ = _0306_ | _0146_;
  assign _0295_ = _0520_ | _0519_;
  assign _0297_ = _0525_ | _0524_;
  assign _0299_ = _0520_ | _0541_;
  assign _0301_ = _0511_ | _0543_;
  assign _0102_ = | { _0520_, _0517_[3], _0517_[1], _0509_ };
  assign _0457_ = _0519_ ? 1'h1 : 1'h0;
  assign _0458_ = _0513_ ? _0003_ : _0000_;
  assign _0460_ = _0509_ ? _0007_ : _0458_;
  assign _0037_ = _0295_ ? _0457_ : _0460_;
  assign _0462_ = _0519_ ? instr_i : { 4'h0, instr_i[8:7], instr_i[12], instr_i[6:2], 8'h12, instr_i[11:9], 9'h023 };
  assign _0464_ = _0513_ ? { 4'h0, instr_i[3:2], instr_i[12], instr_i[6:4], 10'h012, instr_i[11:7], 7'h03 } : { 7'h00, instr_i[6:2], instr_i[11:7], 3'h1, instr_i[11:7], 7'h13 };
  assign _0466_ = _0509_ ? _0035_ : _0464_;
  assign _0031_ = _0295_ ? _0462_ : _0466_;
  assign _0468_ = _0524_ ? instr_i : { 9'h001, instr_i[4:2], 2'h1, instr_i[9:7], 5'h1d, instr_i[9:7], 7'h33 };
  assign _0470_ = _0529_ ? { 9'h001, instr_i[4:2], 2'h1, instr_i[9:7], 5'h11, instr_i[9:7], 7'h33 } : { 9'h081, instr_i[4:2], 2'h1, instr_i[9:7], 5'h01, instr_i[9:7], 7'h33 };
  assign _0472_ = _0527_ ? { 9'h001, instr_i[4:2], 2'h1, instr_i[9:7], 5'h19, instr_i[9:7], 7'h33 } : _0470_;
  assign _0029_ = _0297_ ? _0468_ : _0472_;
  assign _0033_ = _0524_ ? 1'h1 : 1'h0;
  assign _0474_ = _0535_ ? 1'h0 : _0000_;
  assign _0027_ = _0531_ ? _0033_ : _0474_;
  assign _0476_ = _0535_ ? { instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[6:2], 2'h1, instr_i[9:7], 5'h1d, instr_i[9:7], 7'h13 } : { 1'h0, instr_i[10], 5'h00, instr_i[6:2], 2'h1, instr_i[9:7], 5'h15, instr_i[9:7], 7'h13 };
  assign _0025_ = _0531_ ? _0029_ : _0476_;
  assign _0478_ = _0509_ ? _0025_ : _0021_;
  assign _0480_ = _0537_ ? { instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[6:5], instr_i[2], 7'h01, instr_i[9:7], 2'h0, instr_i[13], instr_i[11:10], instr_i[4:3], instr_i[12], 7'h63 } : _0478_;
  assign _0482_ = _0539_ ? { instr_i[12], instr_i[8], instr_i[10:9], instr_i[6], instr_i[7], instr_i[2], instr_i[11], instr_i[5:3], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], 4'h0, _0508_, 7'h6f } : { instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[6:2], instr_i[11:7], 3'h0, instr_i[11:7], 7'h13 };
  assign _0484_ = _0513_ ? { instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[6:2], 8'h00, instr_i[11:7], 7'h13 } : _0482_;
  assign _0017_ = _0102_ ? _0480_ : _0484_;
  assign _0423_ = _0509_ ? _0027_ : _0023_;
  assign _0019_ = _0043_ ? 1'h0 : _0423_;
  assign _0487_ = _0041_ ? 1'h0 : _0015_;
  assign _0011_ = _0541_ ? 1'h1 : _0487_;
  assign _0489_ = _0541_ ? instr_i : { 5'h00, instr_i[5], instr_i[12], 2'h1, instr_i[4:2], 2'h1, instr_i[9:7], 3'h2, instr_i[11:10], instr_i[6], 9'h023 };
  assign _0491_ = _0513_ ? { 5'h00, instr_i[5], instr_i[12:10], instr_i[6], 4'h1, instr_i[9:7], 5'h09, instr_i[4:2], 7'h03 } : { 2'h0, instr_i[10:7], instr_i[12:11], instr_i[5], instr_i[6], 12'h041, instr_i[4:2], 7'h13 };
  assign _0013_ = _0299_ ? _0489_ : _0491_;
  assign _0493_ = _0543_ ? 1'h0 : _0037_;
  assign _0495_ = _0533_ ? _0019_ : _0011_;
  assign illegal_instr_o = _0301_ ? _0493_ : _0495_;
  assign _0497_ = _0543_ ? instr_i : _0031_;
  assign _0499_ = _0533_ ? _0017_ : _0013_;
  assign instr_o = _0301_ ? _0497_ : _0499_;
  assign _0501_ = ! instr_i[12:5];
  assign _0502_ = instr_i[11:7] == 5'h02;
  assign _0504_ = ! { instr_i[12], instr_i[6:2] };
  assign _0505_ = ! instr_i[11:7];
  assign _0506_ = | instr_i[6:2];
  assign is_compressed_o = instr_i[1:0] != 2'h3;
  assign _0508_ = ~ instr_i[15];
  assign _0005_ = _0505_ ? 32'd1048691 : { 12'h000, instr_i[11:7], 15'h00e7 };
  assign _0001_ = _0506_ ? { 7'h00, instr_i[6:2], instr_i[11:7], 3'h0, instr_i[11:7], 7'h33 } : _0005_;
  assign _0039_ = _0506_ ? { 7'h00, instr_i[6:2], 8'h00, instr_i[11:7], 7'h33 } : { 12'h000, instr_i[11:7], 15'h0067 };
  assign _0009_ = _0506_ ? 1'h0 : _0003_;
  assign _0007_ = instr_i[12] ? 1'h0 : _0009_;
  assign _0035_ = instr_i[12] ? _0001_ : _0039_;
  assign _0003_ = _0505_ ? 1'h1 : 1'h0;
  assign _0000_ = instr_i[12] ? 1'h1 : 1'h0;
  assign _0519_ = | _0517_;
  assign _0524_ = | _0522_;
  assign _0522_[0] = { instr_i[12], instr_i[6:5] } == 3'h4;
  assign _0522_[1] = { instr_i[12], instr_i[6:5] } == 3'h5;
  assign _0522_[2] = { instr_i[12], instr_i[6:5] } == 3'h6;
  assign _0522_[3] = { instr_i[12], instr_i[6:5] } == 3'h7;
  assign _0525_ = { instr_i[12], instr_i[6:5] } == 3'h3;
  assign _0527_ = { instr_i[12], instr_i[6:5] } == 3'h2;
  assign _0529_ = { instr_i[12], instr_i[6:5] } == 3'h1;
  assign _0531_ = instr_i[11:10] == 2'h3;
  assign _0535_ = instr_i[11:10] == 2'h2;
  assign _0023_ = _0504_ ? 1'h1 : 1'h0;
  assign _0021_ = _0502_ ? { instr_i[12], instr_i[12], instr_i[12], instr_i[4:3], instr_i[5], instr_i[2], instr_i[6], 24'h010113 } : { instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[6:2], instr_i[11:7], 7'h37 };
  assign _0537_ = | { _0520_, _0517_[3] };
  assign _0539_ = | { _0517_[2], _0517_[0] };
  assign _0015_ = _0501_ ? 1'h1 : 1'h0;
  assign _0541_ = | { _0517_, _0509_ };
  assign _0517_[0] = instr_i[15:13] == 3'h1;
  assign _0517_[1] = instr_i[15:13] == 3'h3;
  assign _0509_ = instr_i[15:13] == 3'h4;
  assign _0517_[2] = instr_i[15:13] == 3'h5;
  assign _0517_[3] = instr_i[15:13] == 3'h7;
  assign _0520_ = instr_i[15:13] == 3'h6;
  assign _0513_ = instr_i[15:13] == 3'h2;
  assign _0515_ = ! instr_i[15:13];
  assign _0533_ = instr_i[1:0] == 2'h1;
  assign _0543_ = instr_i[1:0] == 2'h3;
  assign _0511_ = instr_i[1:0] == 2'h2;
endmodule

module auxy_ibex_load_store_unit(clk_i, rst_ni, data_req_o, data_gnt_i, data_rvalid_i, data_err_i, data_pmp_err_i, data_addr_o, data_we_o, data_be_o, data_wdata_o, data_rdata_i, lsu_we_i, lsu_type_i, lsu_wdata_i, lsu_sign_ext_i, lsu_rdata_o, lsu_rdata_valid_o, lsu_req_i, adder_result_ex_i, addr_incr_req_o
, addr_last_o, lsu_req_done_o, lsu_resp_valid_o, load_err_o, store_err_o, busy_o, perf_load_o, perf_store_o, busy_o_t0, data_req_o_t0, data_we_o_t0, adder_result_ex_i_t0, addr_incr_req_o_t0, addr_last_o_t0, data_addr_o_t0, data_be_o_t0, data_err_i_t0, data_gnt_i_t0, data_pmp_err_i_t0, data_rdata_i_t0, data_rvalid_i_t0
, data_wdata_o_t0, load_err_o_t0, lsu_rdata_o_t0, lsu_rdata_valid_o_t0, lsu_req_done_o_t0, lsu_req_i_t0, lsu_resp_valid_o_t0, lsu_sign_ext_i_t0, lsu_type_i_t0, lsu_wdata_i_t0, lsu_we_i_t0, perf_load_o_t0, perf_store_o_t0, store_err_o_t0);
  wire _0000_;
  wire _0001_;
  wire [3:0] _0002_;
  wire [3:0] _0003_;
  wire _0004_;
  wire _0005_;
  wire _0006_;
  wire [2:0] _0007_;
  wire [2:0] _0008_;
  wire _0009_;
  wire _0010_;
  wire _0011_;
  wire _0012_;
  wire _0013_;
  wire _0014_;
  wire _0015_;
  wire [31:0] _0016_;
  wire [31:0] _0017_;
  wire [31:0] _0018_;
  wire [31:0] _0019_;
  wire _0020_;
  wire _0021_;
  wire _0022_;
  wire [3:0] _0023_;
  wire [3:0] _0024_;
  wire _0025_;
  wire _0026_;
  wire [2:0] _0027_;
  wire [2:0] _0028_;
  wire _0029_;
  wire _0030_;
  wire _0031_;
  wire _0032_;
  wire [31:0] _0033_;
  wire [31:0] _0034_;
  wire [31:0] _0035_;
  wire [31:0] _0036_;
  wire _0037_;
  wire _0038_;
  wire _0039_;
  wire _0040_;
  wire [3:0] _0041_;
  wire [3:0] _0042_;
  wire _0043_;
  wire [2:0] _0044_;
  wire [2:0] _0045_;
  wire _0046_;
  wire _0047_;
  wire _0048_;
  wire _0049_;
  wire [31:0] _0050_;
  wire [31:0] _0051_;
  wire [31:0] _0052_;
  wire [31:0] _0053_;
  wire _0054_;
  wire _0055_;
  wire [3:0] _0056_;
  wire [3:0] _0057_;
  wire _0058_;
  wire _0059_;
  wire [2:0] _0060_;
  wire [2:0] _0061_;
  wire [31:0] _0062_;
  wire [31:0] _0063_;
  wire [31:0] _0064_;
  wire [31:0] _0065_;
  wire _0066_;
  wire _0067_;
  wire [3:0] _0068_;
  wire [3:0] _0069_;
  wire _0070_;
  wire [2:0] _0071_;
  wire [2:0] _0072_;
  wire _0073_;
  wire _0074_;
  wire [3:0] _0075_;
  wire [3:0] _0076_;
  wire _0077_;
  wire [2:0] _0078_;
  wire [2:0] _0079_;
  wire [2:0] _0080_;
  wire [2:0] _0081_;
  wire _0082_;
  wire _0083_;
  wire _0084_;
  wire _0085_;
  wire _0086_;
  wire _0087_;
  wire _0088_;
  wire _0089_;
  wire _0090_;
  wire _0091_;
  wire _0092_;
  wire _0093_;
  wire _0094_;
  wire _0095_;
  wire _0096_;
  wire _0097_;
  wire _0098_;
  wire _0099_;
  wire _0100_;
  wire _0101_;
  wire _0102_;
  wire _0103_;
  wire _0104_;
  wire _0105_;
  wire _0106_;
  wire _0107_;
  wire _0108_;
  wire _0109_;
  wire _0110_;
  wire _0111_;
  wire _0112_;
  wire _0113_;
  wire _0114_;
  wire _0115_;
  wire _0116_;
  wire _0117_;
  wire _0118_;
  wire _0119_;
  wire _0120_;
  wire _0121_;
  wire _0122_;
  wire _0123_;
  wire _0124_;
  wire _0125_;
  wire _0126_;
  wire _0127_;
  wire [2:0] _0128_;
  wire [2:0] _0129_;
  wire [1:0] _0130_;
  wire [1:0] _0131_;
  wire [1:0] _0132_;
  wire [3:0] _0133_;
  wire [1:0] _0134_;
  wire [1:0] _0135_;
  wire [2:0] _0136_;
  wire [1:0] _0137_;
  wire [2:0] _0138_;
  wire [1:0] _0139_;
  wire [2:0] _0140_;
  wire _0141_;
  wire _0142_;
  wire _0143_;
  wire _0144_;
  wire _0145_;
  wire _0146_;
  wire [2:0] _0147_;
  wire [2:0] _0148_;
  wire [2:0] _0149_;
  wire [2:0] _0150_;
  wire [2:0] _0151_;
  wire _0152_;
  wire _0153_;
  wire _0154_;
  wire _0155_;
  wire _0156_;
  wire _0157_;
  wire _0158_;
  wire [31:0] _0159_;
  wire [31:0] _0160_;
  wire [31:0] _0161_;
  wire [31:0] _0162_;
  wire [31:0] _0163_;
  wire [31:0] _0164_;
  wire [31:0] _0165_;
  wire [31:0] _0166_;
  wire [3:0] _0167_;
  wire [3:0] _0168_;
  wire [3:0] _0169_;
  wire [3:0] _0170_;
  wire [3:0] _0171_;
  wire [2:0] _0172_;
  wire _0173_;
  wire _0174_;
  wire _0175_;
  wire _0176_;
  wire _0177_;
  wire [1:0] _0178_;
  wire [2:0] _0179_;
  wire _0180_;
  wire _0181_;
  wire _0182_;
  wire _0183_;
  wire _0184_;
  wire [2:0] _0185_;
  wire [2:0] _0186_;
  wire [2:0] _0187_;
  wire [2:0] _0188_;
  wire [2:0] _0189_;
  wire [1:0] _0190_;
  wire [1:0] _0191_;
  wire [31:0] _0192_;
  wire [1:0] _0193_;
  wire [1:0] _0194_;
  wire [3:0] _0195_;
  wire [1:0] _0196_;
  wire [2:0] _0197_;
  wire _0198_;
  wire _0199_;
  wire _0200_;
  wire _0201_;
  wire _0202_;
  wire _0203_;
  wire _0204_;
  wire _0205_;
  wire _0206_;
  wire _0207_;
  wire _0208_;
  wire _0209_;
  wire _0210_;
  wire _0211_;
  wire _0212_;
  wire _0213_;
  wire _0214_;
  wire _0215_;
  wire _0216_;
  wire _0217_;
  wire _0218_;
  wire _0219_;
  wire _0220_;
  wire _0221_;
  wire _0222_;
  wire _0223_;
  wire _0224_;
  wire _0225_;
  wire _0226_;
  wire _0227_;
  wire _0228_;
  wire _0229_;
  wire _0230_;
  wire _0231_;
  wire _0232_;
  wire _0233_;
  wire _0234_;
  wire _0235_;
  wire _0236_;
  wire _0237_;
  wire _0238_;
  wire _0239_;
  wire _0240_;
  wire _0241_;
  wire _0242_;
  wire _0243_;
  wire _0244_;
  wire _0245_;
  wire _0246_;
  wire _0247_;
  wire _0248_;
  wire _0249_;
  wire _0250_;
  wire _0251_;
  wire _0252_;
  wire _0253_;
  wire _0254_;
  wire _0255_;
  wire _0256_;
  wire _0257_;
  wire _0258_;
  wire _0259_;
  wire _0260_;
  wire _0261_;
  wire _0262_;
  wire _0263_;
  wire _0264_;
  wire _0265_;
  wire _0266_;
  wire _0267_;
  wire _0268_;
  wire [31:0] _0269_;
  wire [31:0] _0270_;
  wire [31:0] _0271_;
  wire [1:0] _0272_;
  wire [1:0] _0273_;
  wire [1:0] _0274_;
  wire [1:0] _0275_;
  wire [1:0] _0276_;
  wire [1:0] _0277_;
  wire _0278_;
  wire _0279_;
  wire _0280_;
  wire _0281_;
  wire _0282_;
  wire _0283_;
  wire _0284_;
  wire _0285_;
  wire _0286_;
  wire _0287_;
  wire _0288_;
  wire _0289_;
  wire [23:0] _0290_;
  wire [23:0] _0291_;
  wire [23:0] _0292_;
  wire _0293_;
  wire _0294_;
  wire _0295_;
  wire [2:0] _0296_;
  wire [2:0] _0297_;
  wire [2:0] _0298_;
  wire [2:0] _0299_;
  wire [1:0] _0300_;
  wire [1:0] _0301_;
  wire [1:0] _0302_;
  wire [1:0] _0303_;
  wire [1:0] _0304_;
  wire [1:0] _0305_;
  wire [3:0] _0306_;
  wire [1:0] _0307_;
  wire [1:0] _0308_;
  wire [1:0] _0309_;
  wire [1:0] _0310_;
  wire [2:0] _0311_;
  wire [1:0] _0312_;
  wire [2:0] _0313_;
  wire [1:0] _0314_;
  wire [2:0] _0315_;
  wire _0316_;
  wire _0317_;
  wire _0318_;
  wire _0319_;
  wire _0320_;
  wire _0321_;
  wire _0322_;
  wire _0323_;
  wire _0324_;
  wire [2:0] _0325_;
  wire [2:0] _0326_;
  wire [2:0] _0327_;
  wire [2:0] _0328_;
  wire [2:0] _0329_;
  wire [2:0] _0330_;
  wire [2:0] _0331_;
  wire [2:0] _0332_;
  wire [2:0] _0333_;
  wire [2:0] _0334_;
  wire [2:0] _0335_;
  wire [2:0] _0336_;
  wire [2:0] _0337_;
  wire [2:0] _0338_;
  wire [2:0] _0339_;
  wire _0340_;
  wire _0341_;
  wire _0342_;
  wire _0343_;
  wire _0344_;
  wire _0345_;
  wire _0346_;
  wire _0347_;
  wire _0348_;
  wire _0349_;
  wire _0350_;
  wire _0351_;
  wire _0352_;
  wire _0353_;
  wire _0354_;
  wire _0355_;
  wire _0356_;
  wire _0357_;
  wire _0358_;
  wire _0359_;
  wire _0360_;
  wire _0361_;
  wire _0362_;
  wire _0363_;
  wire _0364_;
  wire _0365_;
  wire _0366_;
  wire _0367_;
  wire _0368_;
  wire _0369_;
  wire _0370_;
  wire _0371_;
  wire _0372_;
  wire _0373_;
  wire _0374_;
  wire _0375_;
  wire _0376_;
  wire _0377_;
  wire _0378_;
  wire _0379_;
  wire _0380_;
  wire _0381_;
  wire _0382_;
  wire _0383_;
  wire _0384_;
  wire _0385_;
  wire _0386_;
  wire _0387_;
  wire [31:0] _0388_;
  wire [31:0] _0389_;
  wire [31:0] _0390_;
  wire [31:0] _0391_;
  wire [31:0] _0392_;
  wire [31:0] _0393_;
  wire [31:0] _0394_;
  wire [31:0] _0395_;
  wire [31:0] _0396_;
  wire [31:0] _0397_;
  wire [31:0] _0398_;
  wire [31:0] _0399_;
  wire [31:0] _0400_;
  wire [31:0] _0401_;
  wire [31:0] _0402_;
  wire [31:0] _0403_;
  wire [31:0] _0404_;
  wire [31:0] _0405_;
  wire [31:0] _0406_;
  wire [31:0] _0407_;
  wire [31:0] _0408_;
  wire [31:0] _0409_;
  wire [31:0] _0410_;
  wire [31:0] _0411_;
  wire [31:0] _0412_;
  wire [31:0] _0413_;
  wire [31:0] _0414_;
  wire [31:0] _0415_;
  wire [31:0] _0416_;
  wire [31:0] _0417_;
  wire [31:0] _0418_;
  wire [31:0] _0419_;
  wire [31:0] _0420_;
  wire [31:0] _0421_;
  wire [31:0] _0422_;
  wire [31:0] _0423_;
  wire [31:0] _0424_;
  wire [31:0] _0425_;
  wire [31:0] _0426_;
  wire [31:0] _0427_;
  wire [31:0] _0428_;
  wire [31:0] _0429_;
  wire [3:0] _0430_;
  wire [3:0] _0431_;
  wire [3:0] _0432_;
  wire [3:0] _0433_;
  wire [3:0] _0434_;
  wire [3:0] _0435_;
  wire [3:0] _0436_;
  wire [3:0] _0437_;
  wire [3:0] _0438_;
  wire [3:0] _0439_;
  wire [3:0] _0440_;
  wire [3:0] _0441_;
  wire [3:0] _0442_;
  wire [3:0] _0443_;
  wire [3:0] _0444_;
  wire [3:0] _0445_;
  wire [3:0] _0446_;
  wire [3:0] _0447_;
  wire [3:0] _0448_;
  wire [3:0] _0449_;
  wire [3:0] _0450_;
  wire [3:0] _0451_;
  wire [3:0] _0452_;
  wire [3:0] _0453_;
  wire [2:0] _0454_;
  wire _0455_;
  wire _0456_;
  wire _0457_;
  wire _0458_;
  wire _0459_;
  wire _0460_;
  wire _0461_;
  wire _0462_;
  wire _0463_;
  wire _0464_;
  wire _0465_;
  wire _0466_;
  wire _0467_;
  wire _0468_;
  wire _0469_;
  wire [1:0] _0470_;
  wire [2:0] _0471_;
  wire _0472_;
  wire _0473_;
  wire _0474_;
  wire _0475_;
  wire _0476_;
  wire _0477_;
  wire _0478_;
  wire _0479_;
  wire _0480_;
  wire _0481_;
  wire _0482_;
  wire _0483_;
  wire [2:0] _0484_;
  wire [2:0] _0485_;
  wire [2:0] _0486_;
  wire _0487_;
  wire _0488_;
  wire _0489_;
  wire [2:0] _0490_;
  wire [2:0] _0491_;
  wire [2:0] _0492_;
  wire _0493_;
  wire _0494_;
  wire [2:0] _0495_;
  wire [2:0] _0496_;
  wire [2:0] _0497_;
  wire _0498_;
  wire _0499_;
  wire _0500_;
  wire _0501_;
  wire [2:0] _0502_;
  wire [2:0] _0503_;
  wire [2:0] _0504_;
  wire _0505_;
  wire _0506_;
  wire [2:0] _0507_;
  wire [2:0] _0508_;
  wire [2:0] _0509_;
  wire [2:0] _0510_;
  wire [2:0] _0511_;
  wire [2:0] _0512_;
  wire [2:0] _0513_;
  wire _0514_;
  wire _0515_;
  wire _0516_;
  wire _0517_;
  wire _0518_;
  wire _0519_;
  wire _0520_;
  wire _0521_;
  wire _0522_;
  wire _0523_;
  wire _0524_;
  wire [2:0] _0525_;
  wire [2:0] _0526_;
  wire [2:0] _0527_;
  wire [2:0] _0528_;
  wire [1:0] _0529_;
  wire [1:0] _0530_;
  wire [1:0] _0531_;
  wire [1:0] _0532_;
  wire [1:0] _0533_;
  wire [31:0] _0534_;
  wire [31:0] _0535_;
  wire [31:0] _0536_;
  wire [31:0] _0537_;
  wire [31:0] _0538_;
  wire [31:0] _0539_;
  wire [31:0] _0540_;
  wire [31:0] _0541_;
  wire [31:0] _0542_;
  wire [31:0] _0543_;
  wire [31:0] _0544_;
  wire [31:0] _0545_;
  wire [31:0] _0546_;
  wire [31:0] _0547_;
  wire [31:0] _0548_;
  wire [31:0] _0549_;
  wire [31:0] _0550_;
  wire [31:0] _0551_;
  wire [31:0] _0552_;
  wire [31:0] _0553_;
  wire [31:0] _0554_;
  wire [31:0] _0555_;
  wire [31:0] _0556_;
  wire [31:0] _0557_;
  wire [1:0] _0558_;
  wire [1:0] _0559_;
  wire [1:0] _0560_;
  wire [1:0] _0561_;
  wire [1:0] _0562_;
  wire [3:0] _0563_;
  wire [3:0] _0564_;
  wire [3:0] _0565_;
  wire [1:0] _0566_;
  wire [1:0] _0567_;
  wire [1:0] _0568_;
  wire [3:0] _0569_;
  wire [3:0] _0570_;
  wire [3:0] _0571_;
  wire [1:0] _0572_;
  wire [1:0] _0573_;
  wire [1:0] _0574_;
  wire [1:0] _0575_;
  wire [2:0] _0576_;
  wire [2:0] _0577_;
  wire [2:0] _0578_;
  wire [2:0] _0579_;
  wire [2:0] _0580_;
  wire _0581_;
  wire _0582_;
  wire _0583_;
  wire _0584_;
  wire _0585_;
  wire _0586_;
  wire _0587_;
  wire _0588_;
  wire _0589_;
  wire _0590_;
  wire _0591_;
  wire _0592_;
  wire _0593_;
  wire _0594_;
  wire _0595_;
  wire _0596_;
  wire [31:0] _0597_;
  wire [31:0] _0598_;
  wire [31:0] _0599_;
  wire [31:0] _0600_;
  wire [1:0] _0601_;
  wire [1:0] _0602_;
  wire [1:0] _0603_;
  wire [1:0] _0604_;
  wire [1:0] _0605_;
  wire [1:0] _0606_;
  wire [1:0] _0607_;
  wire [1:0] _0608_;
  wire _0609_;
  wire _0610_;
  wire _0611_;
  wire _0612_;
  wire _0613_;
  wire _0614_;
  wire _0615_;
  wire _0616_;
  wire _0617_;
  wire _0618_;
  wire _0619_;
  wire _0620_;
  wire _0621_;
  wire _0622_;
  wire _0623_;
  wire _0624_;
  wire [23:0] _0625_;
  wire [23:0] _0626_;
  wire [23:0] _0627_;
  wire [23:0] _0628_;
  wire _0629_;
  wire _0630_;
  wire _0631_;
  wire _0632_;
  wire [2:0] _0633_;
  wire [1:0] _0634_;
  wire [1:0] _0635_;
  wire [1:0] _0636_;
  wire [5:0] _0637_;
  wire [2:0] _0638_;
  wire [3:0] _0639_;
  wire _0640_;
  wire _0641_;
  wire _0642_;
  wire [2:0] _0643_;
  wire [2:0] _0644_;
  wire [2:0] _0645_;
  wire [2:0] _0646_;
  wire [2:0] _0647_;
  wire [2:0] _0648_;
  wire [2:0] _0649_;
  wire [2:0] _0650_;
  wire [2:0] _0651_;
  wire [2:0] _0652_;
  wire [2:0] _0653_;
  wire [2:0] _0654_;
  wire [2:0] _0655_;
  wire [2:0] _0656_;
  wire [2:0] _0657_;
  wire _0658_;
  wire _0659_;
  wire _0660_;
  wire _0661_;
  wire _0662_;
  wire _0663_;
  wire _0664_;
  wire _0665_;
  wire _0666_;
  wire _0667_;
  wire _0668_;
  wire _0669_;
  wire _0670_;
  wire _0671_;
  wire _0672_;
  wire _0673_;
  wire _0674_;
  wire _0675_;
  wire _0676_;
  wire _0677_;
  wire _0678_;
  wire _0679_;
  wire _0680_;
  wire _0681_;
  wire _0682_;
  wire _0683_;
  wire _0684_;
  wire [31:0] _0685_;
  wire [31:0] _0686_;
  wire [31:0] _0687_;
  wire [31:0] _0688_;
  wire [31:0] _0689_;
  wire [31:0] _0690_;
  wire [31:0] _0691_;
  wire [31:0] _0692_;
  wire [31:0] _0693_;
  wire [31:0] _0694_;
  wire [31:0] _0695_;
  wire [31:0] _0696_;
  wire [31:0] _0697_;
  wire [31:0] _0698_;
  wire [31:0] _0699_;
  wire [31:0] _0700_;
  wire [31:0] _0701_;
  wire [31:0] _0702_;
  wire [31:0] _0703_;
  wire [31:0] _0704_;
  wire [31:0] _0705_;
  wire [31:0] _0706_;
  wire [31:0] _0707_;
  wire [31:0] _0708_;
  wire [31:0] _0709_;
  wire [31:0] _0710_;
  wire [31:0] _0711_;
  wire [31:0] _0712_;
  wire [31:0] _0713_;
  wire [31:0] _0714_;
  wire [3:0] _0715_;
  wire [3:0] _0716_;
  wire [3:0] _0717_;
  wire [3:0] _0718_;
  wire [3:0] _0719_;
  wire [3:0] _0720_;
  wire [3:0] _0721_;
  wire [3:0] _0722_;
  wire [3:0] _0723_;
  wire [3:0] _0724_;
  wire [3:0] _0725_;
  wire [3:0] _0726_;
  wire [3:0] _0727_;
  wire [3:0] _0728_;
  wire [3:0] _0729_;
  wire [3:0] _0730_;
  wire [3:0] _0731_;
  wire _0732_;
  wire _0733_;
  wire _0734_;
  wire _0735_;
  wire _0736_;
  wire _0737_;
  wire _0738_;
  wire _0739_;
  wire _0740_;
  wire [2:0] _0741_;
  wire [2:0] _0742_;
  wire [2:0] _0743_;
  wire _0744_;
  wire _0745_;
  wire [2:0] _0746_;
  wire [2:0] _0747_;
  wire [2:0] _0748_;
  wire _0749_;
  wire [2:0] _0750_;
  wire [2:0] _0751_;
  wire [2:0] _0752_;
  wire _0753_;
  wire [2:0] _0754_;
  wire [2:0] _0755_;
  wire [2:0] _0756_;
  wire [2:0] _0757_;
  wire [2:0] _0758_;
  wire [2:0] _0759_;
  wire [2:0] _0760_;
  wire _0761_;
  wire [31:0] _0762_;
  wire [31:0] _0763_;
  wire [31:0] _0764_;
  wire [31:0] _0765_;
  wire [31:0] _0766_;
  wire [31:0] _0767_;
  wire [31:0] _0768_;
  wire [31:0] _0769_;
  wire [31:0] _0770_;
  wire [31:0] _0771_;
  wire [3:0] _0772_;
  wire [3:0] _0773_;
  wire [3:0] _0774_;
  wire [3:0] _0775_;
  wire [2:0] _0776_;
  wire [2:0] _0777_;
  wire [2:0] _0778_;
  wire [2:0] _0779_;
  wire [31:0] _0780_;
  wire [1:0] _0781_;
  wire [1:0] _0782_;
  wire _0783_;
  wire _0784_;
  wire _0785_;
  wire _0786_;
  wire [23:0] _0787_;
  wire _0788_;
  wire [2:0] _0789_;
  wire [2:0] _0790_;
  wire [2:0] _0791_;
  wire [2:0] _0792_;
  wire _0793_;
  wire _0794_;
  wire _0795_;
  wire _0796_;
  wire _0797_;
  wire _0798_;
  wire _0799_;
  wire _0800_;
  wire _0801_;
  wire _0802_;
  wire _0803_;
  wire _0804_;
  wire [31:0] _0805_;
  wire [31:0] _0806_;
  wire [31:0] _0807_;
  wire [31:0] _0808_;
  wire [31:0] _0809_;
  wire [31:0] _0810_;
  wire [31:0] _0811_;
  wire [31:0] _0812_;
  wire [31:0] _0813_;
  wire [31:0] _0814_;
  wire [31:0] _0815_;
  wire [31:0] _0816_;
  wire [31:0] _0817_;
  wire [31:0] _0818_;
  wire [3:0] _0819_;
  wire [3:0] _0820_;
  wire [3:0] _0821_;
  wire [3:0] _0822_;
  wire [3:0] _0823_;
  wire [3:0] _0824_;
  wire _0825_;
  wire [2:0] _0826_;
  wire _0827_;
  wire [2:0] _0828_;
  wire [2:0] _0829_;
  wire [2:0] _0830_;
  wire [2:0] _0831_;
  wire _0832_;
  wire [31:0] _0833_;
  wire [31:0] _0834_;
  wire [31:0] _0835_;
  wire [31:0] _0836_;
  wire [31:0] _0837_;
  wire [31:0] _0838_;
  wire [31:0] _0839_;
  wire [31:0] _0840_;
  wire [3:0] _0841_;
  wire [3:0] _0842_;
  wire _0843_;
  wire _0844_;
  wire _0845_;
  wire _0846_;
  wire _0847_;
  wire _0848_;
  wire _0849_;
  wire _0850_;
  wire _0851_;
  wire _0852_;
  wire _0853_;
  wire _0854_;
  wire _0855_;
  wire _0856_;
  wire _0857_;
  wire _0858_;
  wire _0859_;
  wire _0860_;
  wire _0861_;
  wire _0862_;
  wire _0863_;
  wire _0864_;
  wire _0865_;
  wire [2:0] _0866_;
  wire [2:0] _0867_;
  wire [2:0] _0868_;
  wire [2:0] _0869_;
  wire [2:0] _0870_;
  wire [2:0] _0871_;
  wire [2:0] _0872_;
  wire [2:0] _0873_;
  wire _0874_;
  wire _0875_;
  wire _0876_;
  wire _0877_;
  wire _0878_;
  wire _0879_;
  wire _0880_;
  wire _0881_;
  wire _0882_;
  wire _0883_;
  wire _0884_;
  wire _0885_;
  wire _0886_;
  wire _0887_;
  wire _0888_;
  wire _0889_;
  wire _0890_;
  wire _0891_;
  wire _0892_;
  wire _0893_;
  wire _0894_;
  wire _0895_;
  wire [31:0] _0896_;
  wire [31:0] _0897_;
  wire [31:0] _0898_;
  wire [31:0] _0899_;
  wire [31:0] _0900_;
  wire [31:0] _0901_;
  wire [31:0] _0902_;
  wire [31:0] _0903_;
  wire [31:0] _0904_;
  wire [31:0] _0905_;
  wire [31:0] _0906_;
  wire [31:0] _0907_;
  wire [31:0] _0908_;
  wire [31:0] _0909_;
  wire [31:0] _0910_;
  wire [31:0] _0911_;
  wire [31:0] _0912_;
  wire [31:0] _0913_;
  wire [3:0] _0914_;
  wire [3:0] _0915_;
  wire [3:0] _0916_;
  wire [3:0] _0917_;
  wire [3:0] _0918_;
  wire [3:0] _0919_;
  wire [3:0] _0920_;
  wire [3:0] _0921_;
  wire [3:0] _0922_;
  wire [3:0] _0923_;
  wire [3:0] _0924_;
  wire [3:0] _0925_;
  wire [3:0] _0926_;
  wire [3:0] _0927_;
  wire _0928_;
  wire _0929_;
  wire _0930_;
  wire _0931_;
  wire _0932_;
  wire _0933_;
  wire _0934_;
  wire _0935_;
  wire _0936_;
  wire _0937_;
  wire _0938_;
  wire _0939_;
  wire _0940_;
  wire _0941_;
  wire _0942_;
  wire _0943_;
  wire _0944_;
  wire _0945_;
  wire _0946_;
  wire _0947_;
  wire _0948_;
  wire _0949_;
  wire _0950_;
  wire _0951_;
  wire _0952_;
  wire _0953_;
  wire _0954_;
  wire _0955_;
  wire _0956_;
  wire _0957_;
  wire [1:0] _0958_;
  wire [1:0] _0959_;
  wire _0960_;
  wire _0961_;
  wire _0962_;
  wire _0963_;
  wire _0964_;
  wire _0965_;
  wire _0966_;
  wire _0967_;
  wire _0968_;
  wire _0969_;
  wire _0970_;
  wire _0971_;
  wire _0972_;
  wire _0973_;
  wire [1:0] _0974_;
  wire [1:0] _0975_;
  wire _0976_;
  wire _0977_;
  wire [2:0] _0978_;
  wire [2:0] _0979_;
  wire [2:0] _0980_;
  wire [2:0] _0981_;
  wire [2:0] _0982_;
  input [31:0] adder_result_ex_i;
  wire [31:0] adder_result_ex_i;
  input [31:0] adder_result_ex_i_t0;
  wire [31:0] adder_result_ex_i_t0;
  output addr_incr_req_o;
  wire addr_incr_req_o;
  output addr_incr_req_o_t0;
  wire addr_incr_req_o_t0;
  output [31:0] addr_last_o;
  reg [31:0] addr_last_o;
  output [31:0] addr_last_o_t0;
  reg [31:0] addr_last_o_t0;
  wire addr_update;
  wire addr_update_t0;
  output busy_o;
  wire busy_o;
  output busy_o_t0;
  wire busy_o_t0;
  input clk_i;
  wire clk_i;
  wire ctrl_update;
  wire ctrl_update_t0;
  output [31:0] data_addr_o;
  wire [31:0] data_addr_o;
  output [31:0] data_addr_o_t0;
  wire [31:0] data_addr_o_t0;
  output [3:0] data_be_o;
  wire [3:0] data_be_o;
  output [3:0] data_be_o_t0;
  wire [3:0] data_be_o_t0;
  input data_err_i;
  wire data_err_i;
  input data_err_i_t0;
  wire data_err_i_t0;
  input data_gnt_i;
  wire data_gnt_i;
  input data_gnt_i_t0;
  wire data_gnt_i_t0;
  wire data_or_pmp_err;
  wire data_or_pmp_err_t0;
  input data_pmp_err_i;
  wire data_pmp_err_i;
  input data_pmp_err_i_t0;
  wire data_pmp_err_i_t0;
  input [31:0] data_rdata_i;
  wire [31:0] data_rdata_i;
  input [31:0] data_rdata_i_t0;
  wire [31:0] data_rdata_i_t0;
  output data_req_o;
  wire data_req_o;
  output data_req_o_t0;
  wire data_req_o_t0;
  input data_rvalid_i;
  wire data_rvalid_i;
  input data_rvalid_i_t0;
  wire data_rvalid_i_t0;
  reg data_sign_ext_q;
  reg data_sign_ext_q_t0;
  reg [1:0] data_type_q;
  reg [1:0] data_type_q_t0;
  output [31:0] data_wdata_o;
  wire [31:0] data_wdata_o;
  output [31:0] data_wdata_o_t0;
  wire [31:0] data_wdata_o_t0;
  output data_we_o;
  wire data_we_o;
  output data_we_o_t0;
  wire data_we_o_t0;
  reg data_we_q;
  reg data_we_q_t0;
  wire handle_misaligned_d;
  wire handle_misaligned_d_t0;
  reg handle_misaligned_q;
  reg handle_misaligned_q_t0;
  output load_err_o;
  wire load_err_o;
  output load_err_o_t0;
  wire load_err_o_t0;
  reg [2:0] ls_fsm_cs;
  reg [2:0] ls_fsm_cs_t0;
  wire [2:0] ls_fsm_ns;
  wire [2:0] ls_fsm_ns_t0;
  wire lsu_err_d;
  wire lsu_err_d_t0;
  reg lsu_err_q;
  reg lsu_err_q_t0;
  output [31:0] lsu_rdata_o;
  wire [31:0] lsu_rdata_o;
  output [31:0] lsu_rdata_o_t0;
  wire [31:0] lsu_rdata_o_t0;
  output lsu_rdata_valid_o;
  wire lsu_rdata_valid_o;
  output lsu_rdata_valid_o_t0;
  wire lsu_rdata_valid_o_t0;
  output lsu_req_done_o;
  wire lsu_req_done_o;
  output lsu_req_done_o_t0;
  wire lsu_req_done_o_t0;
  input lsu_req_i;
  wire lsu_req_i;
  input lsu_req_i_t0;
  wire lsu_req_i_t0;
  output lsu_resp_valid_o;
  wire lsu_resp_valid_o;
  output lsu_resp_valid_o_t0;
  wire lsu_resp_valid_o_t0;
  input lsu_sign_ext_i;
  wire lsu_sign_ext_i;
  input lsu_sign_ext_i_t0;
  wire lsu_sign_ext_i_t0;
  input [1:0] lsu_type_i;
  wire [1:0] lsu_type_i;
  input [1:0] lsu_type_i_t0;
  wire [1:0] lsu_type_i_t0;
  input [31:0] lsu_wdata_i;
  wire [31:0] lsu_wdata_i;
  input [31:0] lsu_wdata_i_t0;
  wire [31:0] lsu_wdata_i_t0;
  input lsu_we_i;
  wire lsu_we_i;
  input lsu_we_i_t0;
  wire lsu_we_i_t0;
  output perf_load_o;
  wire perf_load_o;
  output perf_load_o_t0;
  wire perf_load_o_t0;
  output perf_store_o;
  wire perf_store_o;
  output perf_store_o_t0;
  wire perf_store_o_t0;
  wire pmp_err_d;
  wire pmp_err_d_t0;
  reg pmp_err_q;
  reg pmp_err_q_t0;
  wire [31:0] rdata_b_ext;
  wire [31:0] rdata_b_ext_t0;
  wire [31:0] rdata_h_ext;
  wire [31:0] rdata_h_ext_t0;
  reg [1:0] rdata_offset_q;
  reg [1:0] rdata_offset_q_t0;
  reg [31:8] rdata_q;
  reg [31:8] rdata_q_t0;
  wire rdata_update;
  wire rdata_update_t0;
  wire [31:0] rdata_w_ext;
  wire [31:0] rdata_w_ext_t0;
  input rst_ni;
  wire rst_ni;
  wire split_misaligned_access;
  wire split_misaligned_access_t0;
  output store_err_o;
  wire store_err_o;
  output store_err_o_t0;
  wire store_err_o_t0;
  assign _0082_ = data_gnt_i & _0945_;
  assign lsu_req_done_o = _0949_ & _0934_;
  assign lsu_resp_valid_o = _0953_ & _0936_;
  assign _0084_ = _0936_ & data_rvalid_i;
  assign _0086_ = _0084_ & _0947_;
  assign lsu_rdata_valid_o = _0086_ & _0825_;
  assign _0088_ = data_or_pmp_err & _0825_;
  assign load_err_o = _0088_ & lsu_resp_valid_o;
  assign _0090_ = data_or_pmp_err & data_we_q;
  assign store_err_o = _0090_ & lsu_resp_valid_o;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) ls_fsm_cs_t0 <= 3'h0;
    else ls_fsm_cs_t0 <= ls_fsm_ns_t0;
  assign _0122_ = ~ addr_update;
  assign _0123_ = ~ ctrl_update;
  assign _0124_ = ~ _0110_;
  assign _0125_ = ~ _0112_;
  assign _0126_ = ~ rdata_update;
  assign _0127_ = ~ _0114_;
  assign _0780_ = adder_result_ex_i ^ addr_last_o;
  assign _0781_ = adder_result_ex_i[1:0] ^ rdata_offset_q;
  assign _0782_ = lsu_type_i ^ data_type_q;
  assign _0783_ = lsu_sign_ext_i ^ data_sign_ext_q;
  assign _0784_ = lsu_we_i ^ data_we_q;
  assign _0785_ = handle_misaligned_d ^ handle_misaligned_q;
  assign _0786_ = pmp_err_d ^ pmp_err_q;
  assign _0787_ = data_rdata_i[31:8] ^ rdata_q;
  assign _0788_ = lsu_err_d ^ lsu_err_q;
  assign _0597_ = adder_result_ex_i_t0 | addr_last_o_t0;
  assign _0601_ = adder_result_ex_i_t0[1:0] | rdata_offset_q_t0;
  assign _0605_ = lsu_type_i_t0 | data_type_q_t0;
  assign _0609_ = lsu_sign_ext_i_t0 | data_sign_ext_q_t0;
  assign _0613_ = lsu_we_i_t0 | data_we_q_t0;
  assign _0617_ = handle_misaligned_d_t0 | handle_misaligned_q_t0;
  assign _0621_ = pmp_err_d_t0 | pmp_err_q_t0;
  assign _0625_ = data_rdata_i_t0[31:8] | rdata_q_t0;
  assign _0629_ = lsu_err_d_t0 | lsu_err_q_t0;
  assign _0598_ = _0780_ | _0597_;
  assign _0602_ = _0781_ | _0601_;
  assign _0606_ = _0782_ | _0605_;
  assign _0610_ = _0783_ | _0609_;
  assign _0614_ = _0784_ | _0613_;
  assign _0618_ = _0785_ | _0617_;
  assign _0622_ = _0786_ | _0621_;
  assign _0626_ = _0787_ | _0625_;
  assign _0630_ = _0788_ | _0629_;
  assign _0269_ = { addr_update, addr_update, addr_update, addr_update, addr_update, addr_update, addr_update, addr_update, addr_update, addr_update, addr_update, addr_update, addr_update, addr_update, addr_update, addr_update, addr_update, addr_update, addr_update, addr_update, addr_update, addr_update, addr_update, addr_update, addr_update, addr_update, addr_update, addr_update, addr_update, addr_update, addr_update, addr_update } & adder_result_ex_i_t0;
  assign _0272_ = { ctrl_update, ctrl_update } & adder_result_ex_i_t0[1:0];
  assign _0275_ = { ctrl_update, ctrl_update } & lsu_type_i_t0;
  assign _0278_ = ctrl_update & lsu_sign_ext_i_t0;
  assign _0281_ = ctrl_update & lsu_we_i_t0;
  assign _0284_ = _0110_ & handle_misaligned_d_t0;
  assign _0287_ = _0112_ & pmp_err_d_t0;
  assign _0290_ = { rdata_update, rdata_update, rdata_update, rdata_update, rdata_update, rdata_update, rdata_update, rdata_update, rdata_update, rdata_update, rdata_update, rdata_update, rdata_update, rdata_update, rdata_update, rdata_update, rdata_update, rdata_update, rdata_update, rdata_update, rdata_update, rdata_update, rdata_update, rdata_update } & data_rdata_i_t0[31:8];
  assign _0293_ = _0114_ & lsu_err_d_t0;
  assign _0270_ = { _0122_, _0122_, _0122_, _0122_, _0122_, _0122_, _0122_, _0122_, _0122_, _0122_, _0122_, _0122_, _0122_, _0122_, _0122_, _0122_, _0122_, _0122_, _0122_, _0122_, _0122_, _0122_, _0122_, _0122_, _0122_, _0122_, _0122_, _0122_, _0122_, _0122_, _0122_, _0122_ } & addr_last_o_t0;
  assign _0273_ = { _0123_, _0123_ } & rdata_offset_q_t0;
  assign _0276_ = { _0123_, _0123_ } & data_type_q_t0;
  assign _0279_ = _0123_ & data_sign_ext_q_t0;
  assign _0282_ = _0123_ & data_we_q_t0;
  assign _0285_ = _0124_ & handle_misaligned_q_t0;
  assign _0288_ = _0125_ & pmp_err_q_t0;
  assign _0291_ = { _0126_, _0126_, _0126_, _0126_, _0126_, _0126_, _0126_, _0126_, _0126_, _0126_, _0126_, _0126_, _0126_, _0126_, _0126_, _0126_, _0126_, _0126_, _0126_, _0126_, _0126_, _0126_, _0126_, _0126_ } & rdata_q_t0;
  assign _0294_ = _0127_ & lsu_err_q_t0;
  assign _0271_ = _0598_ & { addr_update_t0, addr_update_t0, addr_update_t0, addr_update_t0, addr_update_t0, addr_update_t0, addr_update_t0, addr_update_t0, addr_update_t0, addr_update_t0, addr_update_t0, addr_update_t0, addr_update_t0, addr_update_t0, addr_update_t0, addr_update_t0, addr_update_t0, addr_update_t0, addr_update_t0, addr_update_t0, addr_update_t0, addr_update_t0, addr_update_t0, addr_update_t0, addr_update_t0, addr_update_t0, addr_update_t0, addr_update_t0, addr_update_t0, addr_update_t0, addr_update_t0, addr_update_t0 };
  assign _0274_ = _0602_ & { ctrl_update_t0, ctrl_update_t0 };
  assign _0277_ = _0606_ & { ctrl_update_t0, ctrl_update_t0 };
  assign _0280_ = _0610_ & ctrl_update_t0;
  assign _0283_ = _0614_ & ctrl_update_t0;
  assign _0286_ = _0618_ & _0111_;
  assign _0289_ = _0622_ & _0113_;
  assign _0292_ = _0626_ & { rdata_update_t0, rdata_update_t0, rdata_update_t0, rdata_update_t0, rdata_update_t0, rdata_update_t0, rdata_update_t0, rdata_update_t0, rdata_update_t0, rdata_update_t0, rdata_update_t0, rdata_update_t0, rdata_update_t0, rdata_update_t0, rdata_update_t0, rdata_update_t0, rdata_update_t0, rdata_update_t0, rdata_update_t0, rdata_update_t0, rdata_update_t0, rdata_update_t0, rdata_update_t0, rdata_update_t0 };
  assign _0295_ = _0630_ & _0115_;
  assign _0599_ = _0269_ | _0270_;
  assign _0603_ = _0272_ | _0273_;
  assign _0607_ = _0275_ | _0276_;
  assign _0611_ = _0278_ | _0279_;
  assign _0615_ = _0281_ | _0282_;
  assign _0619_ = _0284_ | _0285_;
  assign _0623_ = _0287_ | _0288_;
  assign _0627_ = _0290_ | _0291_;
  assign _0631_ = _0293_ | _0294_;
  assign _0600_ = _0599_ | _0271_;
  assign _0604_ = _0603_ | _0274_;
  assign _0608_ = _0607_ | _0277_;
  assign _0612_ = _0611_ | _0280_;
  assign _0616_ = _0615_ | _0283_;
  assign _0620_ = _0619_ | _0286_;
  assign _0624_ = _0623_ | _0289_;
  assign _0628_ = _0627_ | _0292_;
  assign _0632_ = _0631_ | _0295_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) addr_last_o_t0 <= 32'd0;
    else addr_last_o_t0 <= _0600_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) rdata_offset_q_t0 <= 2'h0;
    else rdata_offset_q_t0 <= _0604_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) data_type_q_t0 <= 2'h0;
    else data_type_q_t0 <= _0608_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) data_sign_ext_q_t0 <= 1'h0;
    else data_sign_ext_q_t0 <= _0612_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) data_we_q_t0 <= 1'h0;
    else data_we_q_t0 <= _0616_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) handle_misaligned_q_t0 <= 1'h0;
    else handle_misaligned_q_t0 <= _0620_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) pmp_err_q_t0 <= 1'h0;
    else pmp_err_q_t0 <= _0624_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) rdata_q_t0 <= 24'h000000;
    else rdata_q_t0 <= _0628_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) lsu_err_q_t0 <= 1'h0;
    else lsu_err_q_t0 <= _0632_;
  assign _0241_ = data_gnt_i_t0 & _0945_;
  assign _0244_ = _0950_ & _0934_;
  assign _0247_ = _0633_[1] & _0936_;
  assign _0250_ = busy_o_t0 & data_rvalid_i;
  assign _0253_ = _0085_ & _0947_;
  assign _0256_ = _0087_ & _0825_;
  assign _0259_ = data_or_pmp_err_t0 & _0825_;
  assign _0262_ = _0089_ & lsu_resp_valid_o;
  assign _0265_ = data_or_pmp_err_t0 & data_we_q;
  assign _0266_ = _0091_ & lsu_resp_valid_o;
  assign _0242_ = _0946_ & data_gnt_i;
  assign _0245_ = _0935_ & _0949_;
  assign _0248_ = busy_o_t0 & _0953_;
  assign _0251_ = data_rvalid_i_t0 & _0936_;
  assign _0254_ = data_or_pmp_err_t0 & _0084_;
  assign _0257_ = data_we_q_t0 & _0086_;
  assign _0263_ = lsu_resp_valid_o_t0 & _0088_;
  assign _0260_ = data_we_q_t0 & data_or_pmp_err;
  assign _0267_ = lsu_resp_valid_o_t0 & _0090_;
  assign _0243_ = data_gnt_i_t0 & _0946_;
  assign _0246_ = _0950_ & _0935_;
  assign _0249_ = _0633_[1] & busy_o_t0;
  assign _0252_ = busy_o_t0 & data_rvalid_i_t0;
  assign _0255_ = _0085_ & data_or_pmp_err_t0;
  assign _0258_ = _0087_ & data_we_q_t0;
  assign _0264_ = _0089_ & lsu_resp_valid_o_t0;
  assign _0261_ = data_or_pmp_err_t0 & data_we_q_t0;
  assign _0268_ = _0091_ & lsu_resp_valid_o_t0;
  assign _0587_ = _0241_ | _0242_;
  assign _0588_ = _0244_ | _0245_;
  assign _0589_ = _0247_ | _0248_;
  assign _0590_ = _0250_ | _0251_;
  assign _0591_ = _0253_ | _0254_;
  assign _0592_ = _0256_ | _0257_;
  assign _0593_ = _0259_ | _0260_;
  assign _0594_ = _0262_ | _0263_;
  assign _0595_ = _0265_ | _0260_;
  assign _0596_ = _0266_ | _0267_;
  assign _0083_ = _0587_ | _0243_;
  assign lsu_req_done_o_t0 = _0588_ | _0246_;
  assign lsu_resp_valid_o_t0 = _0589_ | _0249_;
  assign _0085_ = _0590_ | _0252_;
  assign _0087_ = _0591_ | _0255_;
  assign lsu_rdata_valid_o_t0 = _0592_ | _0258_;
  assign _0089_ = _0593_ | _0261_;
  assign load_err_o_t0 = _0594_ | _0264_;
  assign _0091_ = _0595_ | _0261_;
  assign store_err_o_t0 = _0596_ | _0268_;
  assign _0205_ = | { lsu_req_i_t0, data_gnt_i_t0, busy_o_t0 };
  assign _0206_ = | { _0633_[2:1], data_gnt_i_t0 };
  assign _0207_ = | { lsu_req_i_t0, busy_o_t0 };
  assign _0208_ = | { _0040_, _0634_[1] };
  assign _0209_ = | { _0040_, _0635_[1] };
  assign _0211_ = | { _0636_[1], data_rvalid_i_t0 };
  assign _0212_ = | _0633_[2:1];
  assign _0223_ = | ls_fsm_cs_t0;
  assign _0225_ = | data_type_q_t0;
  assign _0226_ = | rdata_offset_q_t0;
  assign _0228_ = | lsu_type_i_t0;
  assign _0128_ = ~ { busy_o_t0, lsu_req_i_t0, data_gnt_i_t0 };
  assign _0129_ = ~ { _0633_[2:1], data_gnt_i_t0 };
  assign _0130_ = ~ { busy_o_t0, lsu_req_i_t0 };
  assign _0131_ = ~ { _0634_[1], _0040_ };
  assign _0132_ = ~ { _0635_[1], _0040_ };
  assign _0134_ = ~ { _0636_[1], data_rvalid_i_t0 };
  assign _0135_ = ~ _0633_[2:1];
  assign _0179_ = ~ ls_fsm_cs_t0;
  assign _0191_ = ~ data_type_q_t0;
  assign _0193_ = ~ rdata_offset_q_t0;
  assign _0178_ = ~ adder_result_ex_i_t0[1:0];
  assign _0196_ = ~ lsu_type_i_t0;
  assign _0296_ = { _0936_, lsu_req_i, data_gnt_i } & _0128_;
  assign _0298_ = { _0956_, _0942_, data_gnt_i } & _0129_;
  assign _0300_ = { _0936_, lsu_req_i } & _0130_;
  assign _0302_ = { _0957_, _0941_ } & _0131_;
  assign _0304_ = { _0955_, _0941_ } & _0132_;
  assign _0307_ = { _0954_, data_rvalid_i } & _0134_;
  assign _0309_ = { _0956_, _0942_ } & _0135_;
  assign _0471_ = ls_fsm_cs & _0179_;
  assign _0530_ = data_type_q & _0191_;
  assign _0558_ = rdata_offset_q & _0193_;
  assign _0470_ = adder_result_ex_i[1:0] & _0178_;
  assign _0572_ = lsu_type_i & _0196_;
  assign _0297_ = 3'h6 & _0128_;
  assign _0299_ = 3'h4 & _0129_;
  assign _0301_ = 2'h2 & _0130_;
  assign _0303_ = 2'h2 & _0131_;
  assign _0305_ = 2'h2 & _0132_;
  assign _0308_ = 2'h2 & _0134_;
  assign _0310_ = 2'h2 & _0135_;
  assign _0525_ = 3'h1 & _0179_;
  assign _0526_ = 3'h4 & _0179_;
  assign _0527_ = 3'h3 & _0179_;
  assign _0528_ = 3'h2 & _0179_;
  assign _0531_ = 2'h2 & _0191_;
  assign _0532_ = 2'h3 & _0191_;
  assign _0533_ = 2'h1 & _0191_;
  assign _0559_ = 2'h3 & _0193_;
  assign _0560_ = 2'h2 & _0193_;
  assign _0561_ = 2'h1 & _0193_;
  assign _0566_ = 2'h3 & _0178_;
  assign _0567_ = 2'h2 & _0178_;
  assign _0568_ = 2'h1 & _0178_;
  assign _0573_ = 2'h2 & _0196_;
  assign _0574_ = 2'h3 & _0196_;
  assign _0575_ = 2'h1 & _0196_;
  assign _0843_ = _0296_ == _0297_;
  assign _0844_ = _0298_ == _0299_;
  assign _0845_ = _0300_ == _0301_;
  assign _0846_ = _0302_ == _0303_;
  assign _0847_ = _0304_ == _0305_;
  assign _0848_ = _0307_ == _0308_;
  assign _0849_ = _0309_ == _0310_;
  assign _0850_ = _0471_ == _0525_;
  assign _0851_ = _0471_ == _0526_;
  assign _0852_ = _0471_ == _0527_;
  assign _0853_ = _0471_ == _0528_;
  assign _0854_ = _0530_ == _0531_;
  assign _0855_ = _0530_ == _0532_;
  assign _0856_ = _0530_ == _0533_;
  assign _0857_ = _0558_ == _0559_;
  assign _0858_ = _0558_ == _0560_;
  assign _0859_ = _0558_ == _0561_;
  assign _0860_ = _0470_ == _0566_;
  assign _0861_ = _0470_ == _0567_;
  assign _0862_ = _0470_ == _0568_;
  assign _0863_ = _0572_ == _0573_;
  assign _0864_ = _0572_ == _0574_;
  assign _0865_ = _0572_ == _0575_;
  assign _0093_ = _0843_ & _0205_;
  assign _0095_ = _0844_ & _0206_;
  assign _0097_ = _0845_ & _0207_;
  assign _0099_ = _0846_ & _0208_;
  assign _0101_ = _0847_ & _0209_;
  assign _0105_ = _0848_ & _0211_;
  assign _0107_ = _0849_ & _0212_;
  assign _0634_[1] = _0850_ & _0223_;
  assign _0636_[1] = _0851_ & _0223_;
  assign _0635_[1] = _0852_ & _0223_;
  assign _0633_[2] = _0853_ & _0223_;
  assign _0959_[0] = _0854_ & _0225_;
  assign _0959_[1] = _0855_ & _0225_;
  assign _0963_ = _0856_ & _0225_;
  assign _0965_ = _0857_ & _0226_;
  assign _0967_ = _0858_ & _0226_;
  assign _0969_ = _0859_ & _0226_;
  assign _0933_ = _0860_ & _0222_;
  assign _0971_ = _0861_ & _0222_;
  assign _0973_ = _0862_ & _0222_;
  assign _0975_[0] = _0863_ & _0228_;
  assign _0975_[1] = _0864_ & _0228_;
  assign _0931_ = _0865_ & _0228_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) addr_last_o <= 32'd0;
    else if (addr_update) addr_last_o <= adder_result_ex_i;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) rdata_offset_q <= 2'h0;
    else if (ctrl_update) rdata_offset_q <= adder_result_ex_i[1:0];
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) data_type_q <= 2'h0;
    else if (ctrl_update) data_type_q <= lsu_type_i;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) data_sign_ext_q <= 1'h0;
    else if (ctrl_update) data_sign_ext_q <= lsu_sign_ext_i;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) data_we_q <= 1'h0;
    else if (ctrl_update) data_we_q <= lsu_we_i;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) handle_misaligned_q <= 1'h0;
    else if (_0110_) handle_misaligned_q <= handle_misaligned_d;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) pmp_err_q <= 1'h0;
    else if (_0112_) pmp_err_q <= pmp_err_d;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) rdata_q <= 24'h000000;
    else if (rdata_update) rdata_q <= data_rdata_i[31:8];
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) lsu_err_q <= 1'h0;
    else if (_0114_) lsu_err_q <= lsu_err_d;
  assign _0455_ = _0929_ & _0943_;
  assign _0458_ = _0931_ & _0932_;
  assign _0456_ = _0944_ & _0928_;
  assign _0459_ = _0933_ & _0930_;
  assign _0457_ = _0929_ & _0944_;
  assign _0460_ = _0931_ & _0933_;
  assign _0732_ = _0455_ | _0456_;
  assign _0733_ = _0458_ | _0459_;
  assign _0938_ = _0732_ | _0457_;
  assign _0940_ = _0733_ | _0460_;
  assign _0210_ = | { _0635_[1], _0634_[1], _0633_[2], busy_o_t0 };
  assign _0213_ = | { _0636_[1], _0633_[2], busy_o_t0 };
  assign _0217_ = | { _0635_[1], _0634_[1] };
  assign _0218_ = | { _0635_[1], _0634_[1], _0633_[2] };
  assign _0219_ = | { _0636_[1], _0633_[2] };
  assign _0220_ = | { _0636_[1], _0635_[1], _0633_[2] };
  assign _0221_ = | ls_fsm_ns_t0;
  assign _0222_ = | adder_result_ex_i_t0[1:0];
  assign _0224_ = | _0959_;
  assign _0227_ = | _0975_;
  assign _0133_ = ~ { _0633_[2], _0635_[1], busy_o_t0, _0634_[1] };
  assign _0136_ = ~ { _0633_[2], _0636_[1], busy_o_t0 };
  assign _0137_ = ~ { _0634_[1], _0635_[1] };
  assign _0138_ = ~ { _0634_[1], _0633_[2], _0635_[1] };
  assign _0139_ = ~ { _0633_[2], _0636_[1] };
  assign _0140_ = ~ { _0633_[2], _0635_[1], _0636_[1] };
  assign _0172_ = ~ ls_fsm_ns_t0;
  assign _0190_ = ~ _0959_;
  assign _0194_ = ~ _0975_;
  assign _0306_ = { _0956_, _0955_, _0936_, _0957_ } & _0133_;
  assign _0311_ = { _0956_, _0954_, _0936_ } & _0136_;
  assign _0312_ = { _0957_, _0955_ } & _0137_;
  assign _0313_ = { _0957_, _0956_, _0955_ } & _0138_;
  assign _0314_ = { _0956_, _0954_ } & _0139_;
  assign _0315_ = { _0956_, _0955_, _0954_ } & _0140_;
  assign _0454_ = ls_fsm_ns & _0172_;
  assign _0529_ = _0958_ & _0190_;
  assign _0562_ = _0974_ & _0194_;
  assign _0229_ = ! _0306_;
  assign _0230_ = ! _0311_;
  assign _0231_ = ! _0312_;
  assign _0232_ = ! _0313_;
  assign _0233_ = ! _0314_;
  assign _0234_ = ! _0315_;
  assign _0235_ = ! _0454_;
  assign _0236_ = ! _0470_;
  assign _0237_ = ! _0471_;
  assign _0238_ = ! _0529_;
  assign _0239_ = ! _0562_;
  assign _0240_ = ! _0572_;
  assign _0103_ = _0229_ & _0210_;
  assign _0109_ = _0230_ & _0213_;
  assign _0117_ = _0231_ & _0217_;
  assign _0121_ = _0232_ & _0218_;
  assign _0119_ = _0233_ & _0219_;
  assign _0204_ = _0234_ & _0220_;
  assign _0935_ = _0235_ & _0221_;
  assign _0944_ = _0236_ & _0222_;
  assign busy_o_t0 = _0237_ & _0223_;
  assign _0961_ = _0238_ & _0224_;
  assign _0977_ = _0239_ & _0227_;
  assign _0929_ = _0240_ & _0228_;
  assign _0173_ = ~ _0937_;
  assign _0174_ = ~ _0939_;
  assign _0461_ = _0938_ & _0174_;
  assign _0467_ = data_gnt_i_t0 & _0176_;
  assign _0462_ = _0940_ & _0173_;
  assign _0468_ = pmp_err_q_t0 & _0177_;
  assign _0463_ = _0938_ & _0940_;
  assign _0469_ = data_gnt_i_t0 & pmp_err_q_t0;
  assign _0734_ = _0461_ | _0462_;
  assign _0736_ = _0467_ | _0468_;
  assign split_misaligned_access_t0 = _0734_ | _0463_;
  assign _0040_ = _0736_ | _0469_;
  assign _0147_ = ~ { _0955_, _0955_, _0955_ };
  assign _0148_ = ~ { _0954_, _0954_, _0954_ };
  assign _0149_ = ~ { _0936_, _0936_, _0936_ };
  assign _0150_ = ~ { _0957_, _0957_, _0957_ };
  assign _0151_ = ~ { _0203_, _0203_, _0203_ };
  assign _0154_ = ~ _0581_;
  assign _0155_ = ~ _0116_;
  assign _0153_ = ~ _0957_;
  assign _0156_ = ~ _0203_;
  assign _0157_ = ~ _0120_;
  assign _0141_ = ~ _0956_;
  assign _0152_ = ~ _0954_;
  assign _0142_ = ~ _0955_;
  assign _0158_ = ~ _0118_;
  assign _0159_ = ~ { _0962_, _0962_, _0962_, _0962_, _0962_, _0962_, _0962_, _0962_, _0962_, _0962_, _0962_, _0962_, _0962_, _0962_, _0962_, _0962_, _0962_, _0962_, _0962_, _0962_, _0962_, _0962_, _0962_, _0962_, _0962_, _0962_, _0962_, _0962_, _0962_, _0962_, _0962_, _0962_ };
  assign _0160_ = ~ { _0960_, _0960_, _0960_, _0960_, _0960_, _0960_, _0960_, _0960_, _0960_, _0960_, _0960_, _0960_, _0960_, _0960_, _0960_, _0960_, _0960_, _0960_, _0960_, _0960_, _0960_, _0960_, _0960_, _0960_, _0960_, _0960_, _0960_, _0960_, _0960_, _0960_, _0960_, _0960_ };
  assign _0161_ = ~ { _0964_, _0964_, _0964_, _0964_, _0964_, _0964_, _0964_, _0964_, _0964_, _0964_, _0964_, _0964_, _0964_, _0964_, _0964_, _0964_, _0964_, _0964_, _0964_, _0964_, _0964_, _0964_, _0964_, _0964_, _0964_, _0964_, _0964_, _0964_, _0964_, _0964_, _0964_, _0964_ };
  assign _0162_ = ~ { _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_ };
  assign _0163_ = ~ { _0583_, _0583_, _0583_, _0583_, _0583_, _0583_, _0583_, _0583_, _0583_, _0583_, _0583_, _0583_, _0583_, _0583_, _0583_, _0583_, _0583_, _0583_, _0583_, _0583_, _0583_, _0583_, _0583_, _0583_, _0583_, _0583_, _0583_, _0583_, _0583_, _0583_, _0583_, _0583_ };
  assign _0164_ = ~ { _0932_, _0932_, _0932_, _0932_, _0932_, _0932_, _0932_, _0932_, _0932_, _0932_, _0932_, _0932_, _0932_, _0932_, _0932_, _0932_, _0932_, _0932_, _0932_, _0932_, _0932_, _0932_, _0932_, _0932_, _0932_, _0932_, _0932_, _0932_, _0932_, _0932_, _0932_, _0932_ };
  assign _0165_ = ~ { _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_ };
  assign _0166_ = ~ { _0585_, _0585_, _0585_, _0585_, _0585_, _0585_, _0585_, _0585_, _0585_, _0585_, _0585_, _0585_, _0585_, _0585_, _0585_, _0585_, _0585_, _0585_, _0585_, _0585_, _0585_, _0585_, _0585_, _0585_, _0585_, _0585_, _0585_, _0585_, _0585_, _0585_, _0585_, _0585_ };
  assign _0167_ = ~ { _0932_, _0932_, _0932_, _0932_ };
  assign _0168_ = ~ { _0972_, _0972_, _0972_, _0972_ };
  assign _0169_ = ~ { _0585_, _0585_, _0585_, _0585_ };
  assign _0170_ = ~ { _0930_, _0930_, _0930_, _0930_ };
  assign _0171_ = ~ { _0976_, _0976_, _0976_, _0976_ };
  assign _0185_ = ~ { data_rvalid_i, data_rvalid_i, data_rvalid_i };
  assign _0175_ = ~ data_rvalid_i;
  assign _0188_ = ~ { _0942_, _0942_, _0942_ };
  assign _0186_ = ~ { _0941_, _0941_, _0941_ };
  assign _0177_ = ~ data_gnt_i;
  assign _0189_ = ~ { lsu_req_i, lsu_req_i, lsu_req_i };
  assign _0181_ = ~ lsu_req_i;
  assign _0192_ = ~ { data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q };
  assign _0195_ = ~ { handle_misaligned_q, handle_misaligned_q, handle_misaligned_q, handle_misaligned_q };
  assign _0197_ = ~ { split_misaligned_access, split_misaligned_access, split_misaligned_access };
  assign _0187_ = ~ { data_gnt_i, data_gnt_i, data_gnt_i };
  assign _0643_ = { _0635_[1], _0635_[1], _0635_[1] } | _0147_;
  assign _0646_ = { _0636_[1], _0636_[1], _0636_[1] } | _0148_;
  assign _0649_ = { busy_o_t0, busy_o_t0, busy_o_t0 } | _0149_;
  assign _0652_ = { _0634_[1], _0634_[1], _0634_[1] } | _0150_;
  assign _0655_ = { _0204_, _0204_, _0204_ } | _0151_;
  assign _0669_ = _0582_ | _0154_;
  assign _0672_ = _0117_ | _0155_;
  assign _0667_ = _0634_[1] | _0153_;
  assign _0679_ = _0204_ | _0156_;
  assign _0682_ = _0121_ | _0157_;
  assign _0658_ = _0633_[2] | _0141_;
  assign _0660_ = _0636_[1] | _0152_;
  assign _0665_ = _0635_[1] | _0142_;
  assign _0684_ = _0119_ | _0158_;
  assign _0685_ = { _0963_, _0963_, _0963_, _0963_, _0963_, _0963_, _0963_, _0963_, _0963_, _0963_, _0963_, _0963_, _0963_, _0963_, _0963_, _0963_, _0963_, _0963_, _0963_, _0963_, _0963_, _0963_, _0963_, _0963_, _0963_, _0963_, _0963_, _0963_, _0963_, _0963_, _0963_, _0963_ } | _0159_;
  assign _0688_ = { _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_ } | _0160_;
  assign _0691_ = { _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_ } | _0161_;
  assign _0694_ = { _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_ } | _0162_;
  assign _0697_ = { _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_ } | _0163_;
  assign _0706_ = { _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_ } | _0164_;
  assign _0709_ = { _0973_, _0973_, _0973_, _0973_, _0973_, _0973_, _0973_, _0973_, _0973_, _0973_, _0973_, _0973_, _0973_, _0973_, _0973_, _0973_, _0973_, _0973_, _0973_, _0973_, _0973_, _0973_, _0973_, _0973_, _0973_, _0973_, _0973_, _0973_, _0973_, _0973_, _0973_, _0973_ } | _0165_;
  assign _0712_ = { _0586_, _0586_, _0586_, _0586_, _0586_, _0586_, _0586_, _0586_, _0586_, _0586_, _0586_, _0586_, _0586_, _0586_, _0586_, _0586_, _0586_, _0586_, _0586_, _0586_, _0586_, _0586_, _0586_, _0586_, _0586_, _0586_, _0586_, _0586_, _0586_, _0586_, _0586_, _0586_ } | _0166_;
  assign _0715_ = { _0933_, _0933_, _0933_, _0933_ } | _0167_;
  assign _0718_ = { _0973_, _0973_, _0973_, _0973_ } | _0168_;
  assign _0721_ = { _0586_, _0586_, _0586_, _0586_ } | _0169_;
  assign _0726_ = { _0931_, _0931_, _0931_, _0931_ } | _0170_;
  assign _0729_ = { _0977_, _0977_, _0977_, _0977_ } | _0171_;
  assign _0741_ = { data_rvalid_i_t0, data_rvalid_i_t0, data_rvalid_i_t0 } | _0185_;
  assign _0754_ = { _0633_[1], _0633_[1], _0633_[1] } | _0188_;
  assign _0746_ = { _0040_, _0040_, _0040_ } | _0186_;
  assign _0758_ = { lsu_req_i_t0, lsu_req_i_t0, lsu_req_i_t0 } | _0189_;
  assign _0762_ = { data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0 } | _0192_;
  assign _0772_ = { handle_misaligned_q_t0, handle_misaligned_q_t0, handle_misaligned_q_t0, handle_misaligned_q_t0 } | _0195_;
  assign _0776_ = { split_misaligned_access_t0, split_misaligned_access_t0, split_misaligned_access_t0 } | _0197_;
  assign _0750_ = { data_gnt_i_t0, data_gnt_i_t0, data_gnt_i_t0 } | _0187_;
  assign _0644_ = { _0635_[1], _0635_[1], _0635_[1] } | { _0955_, _0955_, _0955_ };
  assign _0647_ = { _0636_[1], _0636_[1], _0636_[1] } | { _0954_, _0954_, _0954_ };
  assign _0650_ = { busy_o_t0, busy_o_t0, busy_o_t0 } | { _0936_, _0936_, _0936_ };
  assign _0653_ = { _0634_[1], _0634_[1], _0634_[1] } | { _0957_, _0957_, _0957_ };
  assign _0656_ = { _0204_, _0204_, _0204_ } | { _0203_, _0203_, _0203_ };
  assign _0670_ = _0582_ | _0581_;
  assign _0673_ = _0117_ | _0116_;
  assign _0668_ = _0634_[1] | _0957_;
  assign _0680_ = _0204_ | _0203_;
  assign _0659_ = _0633_[2] | _0956_;
  assign _0661_ = _0636_[1] | _0954_;
  assign _0666_ = _0635_[1] | _0955_;
  assign _0686_ = { _0963_, _0963_, _0963_, _0963_, _0963_, _0963_, _0963_, _0963_, _0963_, _0963_, _0963_, _0963_, _0963_, _0963_, _0963_, _0963_, _0963_, _0963_, _0963_, _0963_, _0963_, _0963_, _0963_, _0963_, _0963_, _0963_, _0963_, _0963_, _0963_, _0963_, _0963_, _0963_ } | { _0962_, _0962_, _0962_, _0962_, _0962_, _0962_, _0962_, _0962_, _0962_, _0962_, _0962_, _0962_, _0962_, _0962_, _0962_, _0962_, _0962_, _0962_, _0962_, _0962_, _0962_, _0962_, _0962_, _0962_, _0962_, _0962_, _0962_, _0962_, _0962_, _0962_, _0962_, _0962_ };
  assign _0689_ = { _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_ } | { _0960_, _0960_, _0960_, _0960_, _0960_, _0960_, _0960_, _0960_, _0960_, _0960_, _0960_, _0960_, _0960_, _0960_, _0960_, _0960_, _0960_, _0960_, _0960_, _0960_, _0960_, _0960_, _0960_, _0960_, _0960_, _0960_, _0960_, _0960_, _0960_, _0960_, _0960_, _0960_ };
  assign _0692_ = { _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_ } | { _0964_, _0964_, _0964_, _0964_, _0964_, _0964_, _0964_, _0964_, _0964_, _0964_, _0964_, _0964_, _0964_, _0964_, _0964_, _0964_, _0964_, _0964_, _0964_, _0964_, _0964_, _0964_, _0964_, _0964_, _0964_, _0964_, _0964_, _0964_, _0964_, _0964_, _0964_, _0964_ };
  assign _0695_ = { _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_ } | { _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_ };
  assign _0698_ = { _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_ } | { _0583_, _0583_, _0583_, _0583_, _0583_, _0583_, _0583_, _0583_, _0583_, _0583_, _0583_, _0583_, _0583_, _0583_, _0583_, _0583_, _0583_, _0583_, _0583_, _0583_, _0583_, _0583_, _0583_, _0583_, _0583_, _0583_, _0583_, _0583_, _0583_, _0583_, _0583_, _0583_ };
  assign _0707_ = { _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_ } | { _0932_, _0932_, _0932_, _0932_, _0932_, _0932_, _0932_, _0932_, _0932_, _0932_, _0932_, _0932_, _0932_, _0932_, _0932_, _0932_, _0932_, _0932_, _0932_, _0932_, _0932_, _0932_, _0932_, _0932_, _0932_, _0932_, _0932_, _0932_, _0932_, _0932_, _0932_, _0932_ };
  assign _0710_ = { _0973_, _0973_, _0973_, _0973_, _0973_, _0973_, _0973_, _0973_, _0973_, _0973_, _0973_, _0973_, _0973_, _0973_, _0973_, _0973_, _0973_, _0973_, _0973_, _0973_, _0973_, _0973_, _0973_, _0973_, _0973_, _0973_, _0973_, _0973_, _0973_, _0973_, _0973_, _0973_ } | { _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_ };
  assign _0713_ = { _0586_, _0586_, _0586_, _0586_, _0586_, _0586_, _0586_, _0586_, _0586_, _0586_, _0586_, _0586_, _0586_, _0586_, _0586_, _0586_, _0586_, _0586_, _0586_, _0586_, _0586_, _0586_, _0586_, _0586_, _0586_, _0586_, _0586_, _0586_, _0586_, _0586_, _0586_, _0586_ } | { _0585_, _0585_, _0585_, _0585_, _0585_, _0585_, _0585_, _0585_, _0585_, _0585_, _0585_, _0585_, _0585_, _0585_, _0585_, _0585_, _0585_, _0585_, _0585_, _0585_, _0585_, _0585_, _0585_, _0585_, _0585_, _0585_, _0585_, _0585_, _0585_, _0585_, _0585_, _0585_ };
  assign _0716_ = { _0933_, _0933_, _0933_, _0933_ } | { _0932_, _0932_, _0932_, _0932_ };
  assign _0719_ = { _0973_, _0973_, _0973_, _0973_ } | { _0972_, _0972_, _0972_, _0972_ };
  assign _0722_ = { _0586_, _0586_, _0586_, _0586_ } | { _0585_, _0585_, _0585_, _0585_ };
  assign _0727_ = { _0931_, _0931_, _0931_, _0931_ } | { _0930_, _0930_, _0930_, _0930_ };
  assign _0730_ = { _0977_, _0977_, _0977_, _0977_ } | { _0976_, _0976_, _0976_, _0976_ };
  assign _0742_ = { data_rvalid_i_t0, data_rvalid_i_t0, data_rvalid_i_t0 } | { data_rvalid_i, data_rvalid_i, data_rvalid_i };
  assign _0744_ = data_rvalid_i_t0 | data_rvalid_i;
  assign _0755_ = { _0633_[1], _0633_[1], _0633_[1] } | { _0942_, _0942_, _0942_ };
  assign _0753_ = _0633_[1] | _0942_;
  assign _0747_ = { _0040_, _0040_, _0040_ } | { _0941_, _0941_, _0941_ };
  assign _0745_ = _0040_ | _0941_;
  assign _0749_ = data_gnt_i_t0 | data_gnt_i;
  assign _0759_ = { lsu_req_i_t0, lsu_req_i_t0, lsu_req_i_t0 } | { lsu_req_i, lsu_req_i, lsu_req_i };
  assign _0761_ = lsu_req_i_t0 | lsu_req_i;
  assign _0677_ = busy_o_t0 | _0936_;
  assign _0763_ = { data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0 } | { data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q };
  assign _0773_ = { handle_misaligned_q_t0, handle_misaligned_q_t0, handle_misaligned_q_t0, handle_misaligned_q_t0 } | { handle_misaligned_q, handle_misaligned_q, handle_misaligned_q, handle_misaligned_q };
  assign _0777_ = { split_misaligned_access_t0, split_misaligned_access_t0, split_misaligned_access_t0 } | { split_misaligned_access, split_misaligned_access, split_misaligned_access };
  assign _0751_ = { data_gnt_i_t0, data_gnt_i_t0, data_gnt_i_t0 } | { data_gnt_i, data_gnt_i, data_gnt_i };
  assign _0325_ = _0061_ & _0643_;
  assign _0328_ = _0867_ & _0646_;
  assign _0331_ = 3'h0 & _0649_;
  assign _0334_ = _0871_ & _0652_;
  assign _0337_ = _0873_ & _0655_;
  assign _0342_ = _0875_ & _0660_;
  assign _0345_ = _0015_ & _0658_;
  assign _0348_ = _0877_ & _0660_;
  assign _0351_ = _0059_ & _0665_;
  assign _0353_ = _0006_ & _0667_;
  assign _0355_ = _0881_ & _0669_;
  assign _0358_ = _0883_ & _0672_;
  assign _0361_ = _0055_ & _0665_;
  assign _0364_ = _0885_ & _0660_;
  assign _0369_ = _0883_ & _0667_;
  assign _0372_ = _0889_ & _0679_;
  assign _0377_ = _0891_ & _0682_;
  assign _0381_ = _0893_ & _0660_;
  assign _0386_ = _0895_ & _0684_;
  assign _0388_ = rdata_w_ext_t0 & _0685_;
  assign _0391_ = _0897_ & _0688_;
  assign _0394_ = _0051_ & _0691_;
  assign _0397_ = _0017_ & _0694_;
  assign _0400_ = _0901_ & _0697_;
  assign _0403_ = _0053_ & _0691_;
  assign _0406_ = _0019_ & _0694_;
  assign _0409_ = _0905_ & _0697_;
  assign _0412_ = { data_rdata_i_t0[15:0], rdata_q_t0[31:16] } & _0691_;
  assign _0415_ = data_rdata_i_t0 & _0694_;
  assign _0418_ = _0909_ & _0697_;
  assign _0421_ = { lsu_wdata_i_t0[15:0], lsu_wdata_i_t0[31:16] } & _0706_;
  assign _0424_ = lsu_wdata_i_t0 & _0709_;
  assign _0427_ = _0913_ & _0712_;
  assign _0436_ = _0917_ & _0721_;
  assign _0440_ = _0921_ & _0721_;
  assign _0430_ = 4'h0 & _0715_;
  assign _0433_ = 4'h0 & _0718_;
  assign _0445_ = _0924_ & _0721_;
  assign _0448_ = _0003_ & _0726_;
  assign _0451_ = _0927_ & _0729_;
  assign _0484_ = ls_fsm_cs_t0 & _0741_;
  assign _0495_ = ls_fsm_cs_t0 & _0750_;
  assign _0502_ = _0072_ & _0754_;
  assign _0490_ = ls_fsm_cs_t0 & _0746_;
  assign _0508_ = _0979_ & _0750_;
  assign _0511_ = ls_fsm_cs_t0 & _0758_;
  assign _0534_ = { 24'h000000, data_rdata_i_t0[31:24] } & _0762_;
  assign _0537_ = { 24'h000000, data_rdata_i_t0[23:16] } & _0762_;
  assign _0540_ = { 24'h000000, data_rdata_i_t0[15:8] } & _0762_;
  assign _0543_ = { 24'h000000, data_rdata_i_t0[7:0] } & _0762_;
  assign _0546_ = { 16'h0000, data_rdata_i_t0[7:0], rdata_q_t0[31:24] } & _0762_;
  assign _0549_ = { 16'h0000, data_rdata_i_t0[31:16] } & _0762_;
  assign _0552_ = { 16'h0000, data_rdata_i_t0[23:8] } & _0762_;
  assign _0555_ = { 16'h0000, data_rdata_i_t0[15:0] } & _0762_;
  assign _0563_ = _0069_ & _0772_;
  assign _0569_ = _0024_ & _0772_;
  assign _0576_ = 3'h0 & _0776_;
  assign _0579_ = 3'h0 & _0750_;
  assign _0326_ = _0079_ & _0644_;
  assign _0329_ = _0081_ & _0647_;
  assign _0332_ = _0008_ & _0650_;
  assign _0335_ = _0045_ & _0653_;
  assign _0338_ = _0869_ & _0656_;
  assign _0340_ = _0030_ & _0659_;
  assign _0343_ = _0047_ & _0661_;
  assign _0346_ = _0032_ & _0659_;
  assign _0349_ = _0049_ & _0661_;
  assign _0356_ = _0879_ & _0670_;
  assign _0359_ = _0040_ & _0673_;
  assign _0362_ = _0067_ & _0666_;
  assign _0365_ = _0074_ & _0661_;
  assign _0367_ = _0001_ & _0677_;
  assign _0370_ = _0040_ & _0668_;
  assign _0373_ = _0887_ & _0680_;
  assign _0375_ = lsu_req_i_t0 & _0677_;
  assign _0379_ = _0021_ & _0659_;
  assign _0382_ = _0038_ & _0661_;
  assign _0384_ = handle_misaligned_q_t0 & _0666_;
  assign _0389_ = rdata_h_ext_t0 & _0686_;
  assign _0392_ = rdata_b_ext_t0 & _0689_;
  assign _0395_ = _0063_ & _0692_;
  assign _0398_ = _0034_ & _0695_;
  assign _0401_ = _0899_ & _0698_;
  assign _0404_ = _0065_ & _0692_;
  assign _0407_ = _0036_ & _0695_;
  assign _0410_ = _0903_ & _0698_;
  assign _0413_ = { data_rdata_i_t0[23:0], rdata_q_t0[31:24] } & _0692_;
  assign _0416_ = { data_rdata_i_t0[7:0], rdata_q_t0 } & _0695_;
  assign _0419_ = _0907_ & _0698_;
  assign _0422_ = { lsu_wdata_i_t0[7:0], lsu_wdata_i_t0[31:8] } & _0707_;
  assign _0425_ = { lsu_wdata_i_t0[23:0], lsu_wdata_i_t0[31:24] } & _0710_;
  assign _0428_ = _0911_ & _0713_;
  assign _0437_ = _0915_ & _0722_;
  assign _0431_ = 4'h0 & _0716_;
  assign _0434_ = 4'h0 & _0719_;
  assign _0441_ = _0919_ & _0722_;
  assign _0449_ = _0057_ & _0727_;
  assign _0452_ = _0076_ & _0730_;
  assign _0485_ = 3'h0 & _0742_;
  assign _0487_ = data_we_q_t0 & _0744_;
  assign _0047_ = data_err_i_t0 & _0744_;
  assign _0049_ = data_pmp_err_i_t0 & _0744_;
  assign _0493_ = lsu_err_q_t0 & _0745_;
  assign _0498_ = data_gnt_i_t0 & _0753_;
  assign _0500_ = _0083_ & _0753_;
  assign _0503_ = _0982_ & _0755_;
  assign _0505_ = data_we_q_t0 & _0753_;
  assign _0030_ = _0946_ & _0753_;
  assign _0032_ = data_pmp_err_i_t0 & _0753_;
  assign _0491_ = 3'h0 & _0747_;
  assign _0509_ = _0979_ & _0751_;
  assign _0026_ = split_misaligned_access_t0 & _0749_;
  assign _0512_ = _0028_ & _0759_;
  assign _0006_ = _0026_ & _0761_;
  assign _0514_ = data_gnt_i_t0 & _0761_;
  assign _0516_ = lsu_we_i_t0 & _0761_;
  assign _0519_ = data_pmp_err_i_t0 & _0761_;
  assign _0521_ = _0013_ & _0677_;
  assign _0523_ = _0011_ & _0677_;
  assign _0535_ = { data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31:24] } & _0763_;
  assign _0538_ = { data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23:16] } & _0763_;
  assign _0541_ = { data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15:8] } & _0763_;
  assign _0544_ = { data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7:0] } & _0763_;
  assign _0547_ = { data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7:0], rdata_q_t0[31:24] } & _0763_;
  assign _0550_ = { data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31:16] } & _0763_;
  assign _0553_ = { data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23:8] } & _0763_;
  assign _0556_ = { data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15:0] } & _0763_;
  assign _0564_ = 4'h0 & _0773_;
  assign _0570_ = _0042_ & _0773_;
  assign _0577_ = 3'h0 & _0777_;
  assign _0496_ = 3'h0 & _0751_;
  assign _0645_ = _0325_ | _0326_;
  assign _0648_ = _0328_ | _0329_;
  assign _0651_ = _0331_ | _0332_;
  assign _0654_ = _0334_ | _0335_;
  assign _0657_ = _0337_ | _0338_;
  assign _0662_ = _0342_ | _0343_;
  assign _0663_ = _0345_ | _0346_;
  assign _0664_ = _0348_ | _0349_;
  assign _0671_ = _0355_ | _0356_;
  assign _0674_ = _0358_ | _0359_;
  assign _0675_ = _0361_ | _0362_;
  assign _0676_ = _0364_ | _0365_;
  assign _0678_ = _0369_ | _0370_;
  assign _0681_ = _0372_ | _0373_;
  assign _0683_ = _0381_ | _0382_;
  assign _0687_ = _0388_ | _0389_;
  assign _0690_ = _0391_ | _0392_;
  assign _0693_ = _0394_ | _0395_;
  assign _0696_ = _0397_ | _0398_;
  assign _0699_ = _0400_ | _0401_;
  assign _0700_ = _0403_ | _0404_;
  assign _0701_ = _0406_ | _0407_;
  assign _0702_ = _0409_ | _0410_;
  assign _0703_ = _0412_ | _0413_;
  assign _0704_ = _0415_ | _0416_;
  assign _0705_ = _0418_ | _0419_;
  assign _0708_ = _0421_ | _0422_;
  assign _0711_ = _0424_ | _0425_;
  assign _0714_ = _0427_ | _0428_;
  assign _0723_ = _0436_ | _0437_;
  assign _0724_ = _0440_ | _0441_;
  assign _0717_ = _0430_ | _0431_;
  assign _0720_ = _0433_ | _0434_;
  assign _0725_ = _0445_ | _0441_;
  assign _0728_ = _0448_ | _0449_;
  assign _0731_ = _0451_ | _0452_;
  assign _0743_ = _0484_ | _0485_;
  assign _0748_ = _0490_ | _0491_;
  assign _0752_ = _0495_ | _0496_;
  assign _0756_ = _0502_ | _0503_;
  assign _0757_ = _0508_ | _0509_;
  assign _0760_ = _0511_ | _0512_;
  assign _0764_ = _0534_ | _0535_;
  assign _0765_ = _0537_ | _0538_;
  assign _0766_ = _0540_ | _0541_;
  assign _0767_ = _0543_ | _0544_;
  assign _0768_ = _0546_ | _0547_;
  assign _0769_ = _0549_ | _0550_;
  assign _0770_ = _0552_ | _0553_;
  assign _0771_ = _0555_ | _0556_;
  assign _0774_ = _0563_ | _0564_;
  assign _0775_ = _0569_ | _0570_;
  assign _0778_ = _0576_ | _0577_;
  assign _0779_ = _0579_ | _0496_;
  assign _0789_ = _0060_ ^ _0078_;
  assign _0790_ = _0866_ ^ _0080_;
  assign _0791_ = _0870_ ^ _0044_;
  assign _0792_ = _0872_ ^ _0868_;
  assign _0793_ = _0009_ ^ _0029_;
  assign _0794_ = _0874_ ^ _0046_;
  assign _0795_ = _0014_ ^ _0031_;
  assign _0796_ = _0876_ ^ _0048_;
  assign _0797_ = _0058_ ^ _0077_;
  assign _0798_ = _0005_ ^ _0043_;
  assign _0799_ = _0880_ ^ _0878_;
  assign _0801_ = _0054_ ^ _0066_;
  assign _0802_ = _0884_ ^ _0073_;
  assign _0800_ = _0882_ ^ _0039_;
  assign _0803_ = _0888_ ^ _0886_;
  assign _0804_ = _0892_ ^ _0037_;
  assign _0805_ = rdata_w_ext ^ rdata_h_ext;
  assign _0806_ = _0896_ ^ rdata_b_ext;
  assign _0807_ = _0050_ ^ _0062_;
  assign _0808_ = _0016_ ^ _0033_;
  assign _0809_ = _0900_ ^ _0898_;
  assign _0810_ = _0052_ ^ _0064_;
  assign _0811_ = _0018_ ^ _0035_;
  assign _0812_ = _0904_ ^ _0902_;
  assign _0813_ = { data_rdata_i[15:0], rdata_q[31:16] } ^ { data_rdata_i[23:0], rdata_q[31:24] };
  assign _0814_ = data_rdata_i ^ { data_rdata_i[7:0], rdata_q };
  assign _0815_ = _0908_ ^ _0906_;
  assign _0816_ = { lsu_wdata_i[15:0], lsu_wdata_i[31:16] } ^ { lsu_wdata_i[7:0], lsu_wdata_i[31:8] };
  assign _0817_ = lsu_wdata_i ^ { lsu_wdata_i[23:0], lsu_wdata_i[31:24] };
  assign _0818_ = _0912_ ^ _0910_;
  assign _0819_ = _0916_ ^ _0914_;
  assign _0820_ = _0920_ ^ _0918_;
  assign _0821_ = _0923_ ^ _0922_;
  assign _0822_ = _0925_ ^ _0918_;
  assign _0823_ = _0002_ ^ _0056_;
  assign _0824_ = _0926_ ^ _0075_;
  assign _0826_ = ls_fsm_cs ^ 3'h4;
  assign _0827_ = _0070_ ^ _0177_;
  assign _0828_ = _0071_ ^ _0981_;
  assign _0829_ = ls_fsm_cs ^ 3'h2;
  assign _0830_ = _0980_ ^ _0978_;
  assign _0831_ = ls_fsm_cs ^ _0027_;
  assign _0833_ = { 24'h000000, data_rdata_i[31:24] } ^ { data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31:24] };
  assign _0834_ = { 24'h000000, data_rdata_i[23:16] } ^ { data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23:16] };
  assign _0835_ = { 24'h000000, data_rdata_i[15:8] } ^ { data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15:8] };
  assign _0836_ = { 24'h000000, data_rdata_i[7:0] } ^ { data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7:0] };
  assign _0837_ = { 16'h0000, data_rdata_i[7:0], rdata_q[31:24] } ^ { data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7:0], rdata_q[31:24] };
  assign _0838_ = { 16'h0000, data_rdata_i[31:16] } ^ { data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31:16] };
  assign _0839_ = { 16'h0000, data_rdata_i[23:8] } ^ { data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23:8] };
  assign _0840_ = { 16'h0000, data_rdata_i[15:0] } ^ { data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15:0] };
  assign _0841_ = _0068_ ^ 4'h1;
  assign _0842_ = _0023_ ^ _0041_;
  assign _0327_ = { _0635_[1], _0635_[1], _0635_[1] } & _0789_;
  assign _0330_ = { _0636_[1], _0636_[1], _0636_[1] } & _0790_;
  assign _0333_ = { busy_o_t0, busy_o_t0, busy_o_t0 } & _0007_;
  assign _0336_ = { _0634_[1], _0634_[1], _0634_[1] } & _0791_;
  assign _0339_ = { _0204_, _0204_, _0204_ } & _0792_;
  assign _0341_ = _0633_[2] & _0793_;
  assign _0344_ = _0636_[1] & _0794_;
  assign _0347_ = _0633_[2] & _0795_;
  assign _0350_ = _0636_[1] & _0796_;
  assign _0352_ = _0635_[1] & _0797_;
  assign _0354_ = _0634_[1] & _0798_;
  assign _0357_ = _0582_ & _0799_;
  assign _0360_ = _0117_ & _0800_;
  assign _0363_ = _0635_[1] & _0801_;
  assign _0366_ = _0636_[1] & _0802_;
  assign _0368_ = busy_o_t0 & _0000_;
  assign _0371_ = _0634_[1] & _0800_;
  assign _0374_ = _0204_ & _0803_;
  assign _0376_ = busy_o_t0 & _0004_;
  assign _0378_ = _0121_ & _0198_;
  assign _0380_ = _0633_[2] & _0020_;
  assign _0383_ = _0636_[1] & _0804_;
  assign _0385_ = _0635_[1] & handle_misaligned_q;
  assign _0387_ = _0119_ & _0199_;
  assign _0390_ = { _0963_, _0963_, _0963_, _0963_, _0963_, _0963_, _0963_, _0963_, _0963_, _0963_, _0963_, _0963_, _0963_, _0963_, _0963_, _0963_, _0963_, _0963_, _0963_, _0963_, _0963_, _0963_, _0963_, _0963_, _0963_, _0963_, _0963_, _0963_, _0963_, _0963_, _0963_, _0963_ } & _0805_;
  assign _0393_ = { _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_ } & _0806_;
  assign _0396_ = { _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_ } & _0807_;
  assign _0399_ = { _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_ } & _0808_;
  assign _0402_ = { _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_ } & _0809_;
  assign _0405_ = { _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_ } & _0810_;
  assign _0408_ = { _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_ } & _0811_;
  assign _0411_ = { _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_ } & _0812_;
  assign _0414_ = { _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_, _0965_ } & _0813_;
  assign _0417_ = { _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_, _0969_ } & _0814_;
  assign _0420_ = { _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_, _0584_ } & _0815_;
  assign _0423_ = { _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_ } & _0816_;
  assign _0426_ = { _0973_, _0973_, _0973_, _0973_, _0973_, _0973_, _0973_, _0973_, _0973_, _0973_, _0973_, _0973_, _0973_, _0973_, _0973_, _0973_, _0973_, _0973_, _0973_, _0973_, _0973_, _0973_, _0973_, _0973_, _0973_, _0973_, _0973_, _0973_, _0973_, _0973_, _0973_, _0973_ } & _0817_;
  assign _0429_ = { _0586_, _0586_, _0586_, _0586_, _0586_, _0586_, _0586_, _0586_, _0586_, _0586_, _0586_, _0586_, _0586_, _0586_, _0586_, _0586_, _0586_, _0586_, _0586_, _0586_, _0586_, _0586_, _0586_, _0586_, _0586_, _0586_, _0586_, _0586_, _0586_, _0586_, _0586_, _0586_ } & _0818_;
  assign _0432_ = { _0933_, _0933_, _0933_, _0933_ } & 4'hc;
  assign _0435_ = { _0973_, _0973_, _0973_, _0973_ } & 4'h3;
  assign _0438_ = { _0586_, _0586_, _0586_, _0586_ } & _0819_;
  assign _0439_ = { _0973_, _0973_, _0973_, _0973_ } & 4'h5;
  assign _0442_ = { _0586_, _0586_, _0586_, _0586_ } & _0820_;
  assign _0446_ = { _0586_, _0586_, _0586_, _0586_ } & _0821_;
  assign _0443_ = { _0933_, _0933_, _0933_, _0933_ } & 4'h4;
  assign _0444_ = { _0973_, _0973_, _0973_, _0973_ } & 4'h1;
  assign _0447_ = { _0586_, _0586_, _0586_, _0586_ } & _0822_;
  assign _0450_ = { _0931_, _0931_, _0931_, _0931_ } & _0823_;
  assign _0453_ = { _0977_, _0977_, _0977_, _0977_ } & _0824_;
  assign _0486_ = { data_rvalid_i_t0, data_rvalid_i_t0, data_rvalid_i_t0 } & ls_fsm_cs;
  assign _0488_ = data_rvalid_i_t0 & _0825_;
  assign _0489_ = data_rvalid_i_t0 & _0180_;
  assign _0492_ = { _0040_, _0040_, _0040_ } & ls_fsm_cs;
  assign _0494_ = _0040_ & _0183_;
  assign _0497_ = { data_gnt_i_t0, data_gnt_i_t0, data_gnt_i_t0 } & _0826_;
  assign _0499_ = _0633_[1] & _0827_;
  assign _0501_ = _0633_[1] & _0082_;
  assign _0504_ = { _0633_[1], _0633_[1], _0633_[1] } & _0828_;
  assign _0506_ = _0633_[1] & _0825_;
  assign _0507_ = { _0040_, _0040_, _0040_ } & _0829_;
  assign _0510_ = { data_gnt_i_t0, data_gnt_i_t0, data_gnt_i_t0 } & _0830_;
  assign _0513_ = { lsu_req_i_t0, lsu_req_i_t0, lsu_req_i_t0 } & _0831_;
  assign _0515_ = lsu_req_i_t0 & _0022_;
  assign _0517_ = lsu_req_i_t0 & lsu_we_i;
  assign _0518_ = lsu_req_i_t0 & _0832_;
  assign _0520_ = lsu_req_i_t0 & data_pmp_err_i;
  assign _0522_ = busy_o_t0 & _0012_;
  assign _0524_ = busy_o_t0 & _0010_;
  assign _0536_ = { data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0 } & _0833_;
  assign _0539_ = { data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0 } & _0834_;
  assign _0542_ = { data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0 } & _0835_;
  assign _0545_ = { data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0 } & _0836_;
  assign _0548_ = { data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0 } & _0837_;
  assign _0551_ = { data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0 } & _0838_;
  assign _0554_ = { data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0 } & _0839_;
  assign _0557_ = { data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0 } & _0840_;
  assign _0565_ = { handle_misaligned_q_t0, handle_misaligned_q_t0, handle_misaligned_q_t0, handle_misaligned_q_t0 } & _0841_;
  assign _0571_ = { handle_misaligned_q_t0, handle_misaligned_q_t0, handle_misaligned_q_t0, handle_misaligned_q_t0 } & _0842_;
  assign _0578_ = { split_misaligned_access_t0, split_misaligned_access_t0, split_misaligned_access_t0 } & 3'h2;
  assign _0580_ = { data_gnt_i_t0, data_gnt_i_t0, data_gnt_i_t0 } & 3'h3;
  assign _0867_ = _0327_ | _0645_;
  assign _0869_ = _0330_ | _0648_;
  assign _0871_ = _0333_ | _0651_;
  assign _0873_ = _0336_ | _0654_;
  assign ls_fsm_ns_t0 = _0339_ | _0657_;
  assign _0875_ = _0341_ | _0340_;
  assign lsu_err_d_t0 = _0344_ | _0662_;
  assign _0877_ = _0347_ | _0663_;
  assign pmp_err_d_t0 = _0350_ | _0664_;
  assign _0879_ = _0352_ | _0351_;
  assign _0881_ = _0354_ | _0353_;
  assign handle_misaligned_d_t0 = _0357_ | _0671_;
  assign ctrl_update_t0 = _0360_ | _0674_;
  assign _0885_ = _0363_ | _0675_;
  assign _0887_ = _0366_ | _0676_;
  assign _0883_ = _0368_ | _0367_;
  assign _0889_ = _0371_ | _0678_;
  assign addr_update_t0 = _0374_ | _0681_;
  assign _0891_ = _0376_ | _0375_;
  assign data_req_o_t0 = _0378_ | _0377_;
  assign _0893_ = _0380_ | _0379_;
  assign rdata_update_t0 = _0383_ | _0683_;
  assign _0895_ = _0385_ | _0384_;
  assign addr_incr_req_o_t0 = _0387_ | _0386_;
  assign _0897_ = _0390_ | _0687_;
  assign lsu_rdata_o_t0 = _0393_ | _0690_;
  assign _0899_ = _0396_ | _0693_;
  assign _0901_ = _0399_ | _0696_;
  assign rdata_b_ext_t0 = _0402_ | _0699_;
  assign _0903_ = _0405_ | _0700_;
  assign _0905_ = _0408_ | _0701_;
  assign rdata_h_ext_t0 = _0411_ | _0702_;
  assign _0907_ = _0414_ | _0703_;
  assign _0909_ = _0417_ | _0704_;
  assign rdata_w_ext_t0 = _0420_ | _0705_;
  assign _0911_ = _0423_ | _0708_;
  assign _0913_ = _0426_ | _0711_;
  assign data_wdata_o_t0 = _0429_ | _0714_;
  assign _0915_ = _0432_ | _0717_;
  assign _0917_ = _0435_ | _0720_;
  assign _0076_ = _0438_ | _0723_;
  assign _0921_ = _0439_ | _0720_;
  assign _0069_ = _0442_ | _0724_;
  assign _0042_ = _0446_ | _0725_;
  assign _0919_ = _0443_ | _0717_;
  assign _0924_ = _0444_ | _0720_;
  assign _0024_ = _0447_ | _0725_;
  assign _0927_ = _0450_ | _0728_;
  assign data_be_o_t0 = _0453_ | _0731_;
  assign _0081_ = _0486_ | _0743_;
  assign _0038_ = _0488_ | _0487_;
  assign _0074_ = _0489_ | _0047_;
  assign _0079_ = _0492_ | _0748_;
  assign _0067_ = _0494_ | _0493_;
  assign _0072_ = _0497_ | _0752_;
  assign _0059_ = _0499_ | _0498_;
  assign _0055_ = _0501_ | _0500_;
  assign _0061_ = _0504_ | _0756_;
  assign _0021_ = _0506_ | _0505_;
  assign _0045_ = _0507_ | _0748_;
  assign _0028_ = _0510_ | _0757_;
  assign _0008_ = _0513_ | _0760_;
  assign _0001_ = _0515_ | _0514_;
  assign _0013_ = _0517_ | _0516_;
  assign _0011_ = _0518_ | _0516_;
  assign _0015_ = _0520_ | _0519_;
  assign perf_store_o_t0 = _0522_ | _0521_;
  assign perf_load_o_t0 = _0524_ | _0523_;
  assign _0063_ = _0536_ | _0764_;
  assign _0051_ = _0539_ | _0765_;
  assign _0034_ = _0542_ | _0766_;
  assign _0017_ = _0545_ | _0767_;
  assign _0065_ = _0548_ | _0768_;
  assign _0053_ = _0551_ | _0769_;
  assign _0036_ = _0554_ | _0770_;
  assign _0019_ = _0557_ | _0771_;
  assign _0057_ = _0565_ | _0774_;
  assign _0003_ = _0571_ | _0775_;
  assign _0979_ = _0578_ | _0778_;
  assign _0982_ = _0580_ | _0779_;
  assign _0092_ = { _0936_, lsu_req_i, data_gnt_i } != 3'h6;
  assign _0094_ = { _0956_, _0942_, data_gnt_i } != 3'h4;
  assign _0096_ = { _0936_, lsu_req_i } != 2'h2;
  assign _0098_ = { _0957_, _0941_ } != 2'h2;
  assign _0100_ = { _0955_, _0941_ } != 2'h2;
  assign _0102_ = | { _0956_, _0955_, _0936_, _0957_ };
  assign _0104_ = { _0954_, data_rvalid_i } != 2'h2;
  assign _0106_ = { _0956_, _0942_ } != 2'h2;
  assign _0108_ = | { _0956_, _0954_, _0936_ };
  assign _0110_ = & { _0098_, _0102_, _0100_, _0094_, _0092_, _0096_ };
  assign _0112_ = & { _0108_, _0106_, _0104_ };
  assign _0114_ = & { _0108_, _0106_, _0104_, _0096_ };
  assign _0198_ = ~ _0890_;
  assign _0199_ = ~ _0894_;
  assign _0116_ = | { _0957_, _0955_ };
  assign _0120_ = | { _0957_, _0956_, _0955_ };
  assign _0143_ = ~ _0966_;
  assign _0145_ = ~ _0970_;
  assign _0183_ = ~ lsu_err_q;
  assign _0184_ = ~ _0951_;
  assign _0144_ = ~ _0964_;
  assign _0146_ = ~ _0932_;
  assign _0182_ = ~ busy_o;
  assign _0180_ = ~ data_err_i;
  assign _0176_ = ~ pmp_err_q;
  assign _0316_ = _0633_[2] & _0142_;
  assign _0319_ = _0967_ & _0144_;
  assign _0322_ = _0971_ & _0146_;
  assign _0472_ = data_err_i_t0 & _0176_;
  assign _0475_ = lsu_req_i_t0 & _0182_;
  assign _0478_ = lsu_err_q_t0 & _0180_;
  assign _0481_ = _0952_ & _0176_;
  assign _0464_ = data_rvalid_i_t0 & _0176_;
  assign _0317_ = _0635_[1] & _0141_;
  assign _0320_ = _0965_ & _0143_;
  assign _0323_ = _0933_ & _0145_;
  assign _0473_ = pmp_err_q_t0 & _0180_;
  assign _0476_ = busy_o_t0 & _0181_;
  assign _0479_ = data_err_i_t0 & _0183_;
  assign _0482_ = pmp_err_q_t0 & _0184_;
  assign _0465_ = pmp_err_q_t0 & _0175_;
  assign _0318_ = _0633_[2] & _0635_[1];
  assign _0321_ = _0967_ & _0965_;
  assign _0324_ = _0971_ & _0933_;
  assign _0474_ = data_err_i_t0 & pmp_err_q_t0;
  assign _0477_ = lsu_req_i_t0 & busy_o_t0;
  assign _0480_ = lsu_err_q_t0 & data_err_i_t0;
  assign _0483_ = _0952_ & pmp_err_q_t0;
  assign _0466_ = data_rvalid_i_t0 & pmp_err_q_t0;
  assign _0640_ = _0316_ | _0317_;
  assign _0641_ = _0319_ | _0320_;
  assign _0642_ = _0322_ | _0323_;
  assign _0737_ = _0472_ | _0473_;
  assign _0738_ = _0475_ | _0476_;
  assign _0739_ = _0478_ | _0479_;
  assign _0740_ = _0481_ | _0482_;
  assign _0735_ = _0464_ | _0465_;
  assign _0582_ = _0640_ | _0318_;
  assign _0584_ = _0641_ | _0321_;
  assign _0586_ = _0642_ | _0324_;
  assign _0946_ = _0737_ | _0474_;
  assign _0950_ = _0738_ | _0477_;
  assign _0952_ = _0739_ | _0480_;
  assign data_or_pmp_err_t0 = _0740_ | _0483_;
  assign _0633_[1] = _0735_ | _0466_;
  assign _0118_ = | { _0956_, _0954_ };
  assign _0203_ = | { _0956_, _0955_, _0954_ };
  assign _0581_ = _0956_ | _0955_;
  assign _0583_ = _0966_ | _0964_;
  assign _0585_ = _0970_ | _0932_;
  assign _0866_ = _0955_ ? _0078_ : _0060_;
  assign _0868_ = _0954_ ? _0080_ : _0866_;
  assign _0870_ = _0936_ ? _0007_ : 3'h0;
  assign _0872_ = _0957_ ? _0044_ : _0870_;
  assign ls_fsm_ns = _0203_ ? _0868_ : _0872_;
  assign _0874_ = _0956_ ? _0029_ : _0009_;
  assign lsu_err_d = _0954_ ? _0046_ : _0874_;
  assign _0876_ = _0956_ ? _0031_ : _0014_;
  assign pmp_err_d = _0954_ ? _0048_ : _0876_;
  assign _0878_ = _0955_ ? _0077_ : _0058_;
  assign _0880_ = _0957_ ? _0043_ : _0005_;
  assign handle_misaligned_d = _0581_ ? _0878_ : _0880_;
  assign ctrl_update = _0116_ ? _0039_ : _0882_;
  assign _0884_ = _0955_ ? _0066_ : _0054_;
  assign _0886_ = _0954_ ? _0073_ : _0884_;
  assign _0882_ = _0936_ ? _0000_ : 1'h0;
  assign _0888_ = _0957_ ? _0039_ : _0882_;
  assign addr_update = _0203_ ? _0886_ : _0888_;
  assign _0890_ = _0936_ ? _0004_ : 1'h0;
  assign data_req_o = _0120_ ? 1'h1 : _0890_;
  assign _0892_ = _0956_ ? _0020_ : 1'h0;
  assign rdata_update = _0954_ ? _0037_ : _0892_;
  assign _0894_ = _0955_ ? handle_misaligned_q : 1'h0;
  assign addr_incr_req_o = _0118_ ? 1'h1 : _0894_;
  assign _0896_ = _0962_ ? rdata_h_ext : rdata_w_ext;
  assign lsu_rdata_o = _0960_ ? rdata_b_ext : _0896_;
  assign _0898_ = _0964_ ? _0062_ : _0050_;
  assign _0900_ = _0968_ ? _0033_ : _0016_;
  assign rdata_b_ext = _0583_ ? _0898_ : _0900_;
  assign _0902_ = _0964_ ? _0064_ : _0052_;
  assign _0904_ = _0968_ ? _0035_ : _0018_;
  assign rdata_h_ext = _0583_ ? _0902_ : _0904_;
  assign _0906_ = _0964_ ? { data_rdata_i[23:0], rdata_q[31:24] } : { data_rdata_i[15:0], rdata_q[31:16] };
  assign _0908_ = _0968_ ? { data_rdata_i[7:0], rdata_q } : data_rdata_i;
  assign rdata_w_ext = _0583_ ? _0906_ : _0908_;
  assign _0910_ = _0932_ ? { lsu_wdata_i[7:0], lsu_wdata_i[31:8] } : { lsu_wdata_i[15:0], lsu_wdata_i[31:16] };
  assign _0912_ = _0972_ ? { lsu_wdata_i[23:0], lsu_wdata_i[31:24] } : lsu_wdata_i;
  assign data_wdata_o = _0585_ ? _0910_ : _0912_;
  assign _0914_ = _0932_ ? 4'h8 : 4'h4;
  assign _0916_ = _0972_ ? 4'h2 : 4'h1;
  assign _0075_ = _0585_ ? _0914_ : _0916_;
  assign _0920_ = _0972_ ? 4'h6 : 4'h3;
  assign _0068_ = _0585_ ? _0918_ : _0920_;
  assign _0922_ = _0932_ ? 4'h7 : 4'h3;
  assign _0923_ = _0972_ ? 4'h1 : 4'h0;
  assign _0041_ = _0585_ ? _0922_ : _0923_;
  assign _0918_ = _0932_ ? 4'h8 : 4'hc;
  assign _0925_ = _0972_ ? 4'he : 4'hf;
  assign _0023_ = _0585_ ? _0918_ : _0925_;
  assign _0926_ = _0930_ ? _0056_ : _0002_;
  assign data_be_o = _0976_ ? _0075_ : _0926_;
  assign _0214_ = | { _0103_, _0101_, _0099_, _0097_, _0095_, _0093_ };
  assign _0215_ = | { _0109_, _0107_, _0105_ };
  assign _0216_ = | { _0109_, _0107_, _0105_, _0097_ };
  assign _0637_ = { _0098_, _0102_, _0100_, _0094_, _0092_, _0096_ } | { _0099_, _0103_, _0101_, _0095_, _0093_, _0097_ };
  assign _0638_ = { _0108_, _0106_, _0104_ } | { _0109_, _0107_, _0105_ };
  assign _0639_ = { _0108_, _0106_, _0104_, _0096_ } | { _0109_, _0107_, _0105_, _0097_ };
  assign _0200_ = & _0637_;
  assign _0201_ = & _0638_;
  assign _0202_ = & _0639_;
  assign _0111_ = _0214_ & _0200_;
  assign _0113_ = _0215_ & _0201_;
  assign _0115_ = _0216_ & _0202_;
  assign _0934_ = ! ls_fsm_ns;
  assign _0937_ = _0928_ && _0943_;
  assign _0939_ = _0930_ && _0932_;
  assign split_misaligned_access = _0937_ || _0939_;
  assign _0942_ = data_rvalid_i || pmp_err_q;
  assign _0941_ = data_gnt_i || pmp_err_q;
  assign _0943_ = | adder_result_ex_i[1:0];
  assign busy_o = | ls_fsm_cs;
  assign _0832_ = ~ lsu_we_i;
  assign _0945_ = ~ _0948_;
  assign _0947_ = ~ data_or_pmp_err;
  assign _0825_ = ~ data_we_q;
  assign _0948_ = data_err_i | pmp_err_q;
  assign _0949_ = lsu_req_i | busy_o;
  assign _0951_ = lsu_err_q | data_err_i;
  assign data_or_pmp_err = _0951_ | pmp_err_q;
  assign _0953_ = data_rvalid_i | pmp_err_q;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) ls_fsm_cs <= 3'h0;
    else ls_fsm_cs <= ls_fsm_ns;
  assign _0080_ = data_rvalid_i ? 3'h0 : ls_fsm_cs;
  assign _0037_ = data_rvalid_i ? _0825_ : 1'h0;
  assign _0073_ = data_rvalid_i ? _0180_ : 1'h0;
  assign _0046_ = data_rvalid_i ? data_err_i : 1'hx;
  assign _0048_ = data_rvalid_i ? data_pmp_err_i : 1'hx;
  assign _0077_ = _0941_ ? 1'h0 : 1'hx;
  assign _0078_ = _0941_ ? 3'h0 : ls_fsm_cs;
  assign _0066_ = _0941_ ? _0183_ : 1'h0;
  assign _0070_ = data_gnt_i ? 1'h0 : 1'hx;
  assign _0071_ = data_gnt_i ? 3'h4 : ls_fsm_cs;
  assign _0058_ = _0942_ ? _0177_ : _0070_;
  assign _0054_ = _0942_ ? _0082_ : 1'h0;
  assign _0060_ = _0942_ ? _0981_ : _0071_;
  assign _0020_ = _0942_ ? _0825_ : 1'h0;
  assign _0029_ = _0942_ ? _0948_ : 1'hx;
  assign _0031_ = _0942_ ? data_pmp_err_i : 1'hx;
  assign _0044_ = _0941_ ? 3'h2 : ls_fsm_cs;
  assign _0043_ = _0941_ ? 1'h1 : 1'hx;
  assign _0039_ = _0941_ ? 1'h1 : 1'h0;
  assign _0027_ = data_gnt_i ? _0978_ : _0980_;
  assign _0025_ = data_gnt_i ? split_misaligned_access : 1'hx;
  assign _0022_ = data_gnt_i ? 1'h1 : 1'h0;
  assign _0007_ = lsu_req_i ? _0027_ : ls_fsm_cs;
  assign _0005_ = lsu_req_i ? _0025_ : 1'hx;
  assign _0000_ = lsu_req_i ? _0022_ : 1'h0;
  assign _0012_ = lsu_req_i ? lsu_we_i : 1'h0;
  assign _0010_ = lsu_req_i ? _0832_ : 1'h0;
  assign _0009_ = lsu_req_i ? 1'h0 : 1'hx;
  assign _0014_ = lsu_req_i ? data_pmp_err_i : 1'h0;
  assign _0004_ = lsu_req_i ? 1'h1 : 1'h0;
  assign perf_store_o = _0936_ ? _0012_ : 1'h0;
  assign perf_load_o = _0936_ ? _0010_ : 1'h0;
  assign _0957_ = ls_fsm_cs == 3'h1;
  assign _0936_ = ! ls_fsm_cs;
  assign _0954_ = ls_fsm_cs == 3'h4;
  assign _0955_ = ls_fsm_cs == 3'h3;
  assign _0956_ = ls_fsm_cs == 3'h2;
  assign _0960_ = | _0958_;
  assign _0958_[0] = data_type_q == 2'h2;
  assign _0958_[1] = data_type_q == 2'h3;
  assign _0962_ = data_type_q == 2'h1;
  assign _0062_ = data_sign_ext_q ? { data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31:24] } : { 24'h000000, data_rdata_i[31:24] };
  assign _0050_ = data_sign_ext_q ? { data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23:16] } : { 24'h000000, data_rdata_i[23:16] };
  assign _0033_ = data_sign_ext_q ? { data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15:8] } : { 24'h000000, data_rdata_i[15:8] };
  assign _0016_ = data_sign_ext_q ? { data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7:0] } : { 24'h000000, data_rdata_i[7:0] };
  assign _0064_ = data_sign_ext_q ? { data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7:0], rdata_q[31:24] } : { 16'h0000, data_rdata_i[7:0], rdata_q[31:24] };
  assign _0052_ = data_sign_ext_q ? { data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31:16] } : { 16'h0000, data_rdata_i[31:16] };
  assign _0035_ = data_sign_ext_q ? { data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23:8] } : { 16'h0000, data_rdata_i[23:8] };
  assign _0018_ = data_sign_ext_q ? { data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15:0] } : { 16'h0000, data_rdata_i[15:0] };
  assign _0964_ = rdata_offset_q == 2'h3;
  assign _0966_ = rdata_offset_q == 2'h2;
  assign _0968_ = rdata_offset_q == 2'h1;
  assign _0976_ = | _0974_;
  assign _0056_ = handle_misaligned_q ? 4'h1 : _0068_;
  assign _0932_ = adder_result_ex_i[1:0] == 2'h3;
  assign _0970_ = adder_result_ex_i[1:0] == 2'h2;
  assign _0972_ = adder_result_ex_i[1:0] == 2'h1;
  assign _0002_ = handle_misaligned_q ? _0041_ : _0023_;
  assign _0974_[0] = lsu_type_i == 2'h2;
  assign _0974_[1] = lsu_type_i == 2'h3;
  assign _0930_ = lsu_type_i == 2'h1;
  assign _0928_ = ! lsu_type_i;
  assign _0978_ = split_misaligned_access ? 3'h2 : 3'h0;
  assign _0980_ = split_misaligned_access ? 3'h1 : 3'h3;
  assign _0981_ = data_gnt_i ? 3'h0 : 3'h3;
  assign _0633_[0] = data_gnt_i_t0;
  assign _0634_[0] = _0040_;
  assign _0635_[0] = _0040_;
  assign _0636_[0] = data_rvalid_i_t0;
  assign data_addr_o = { adder_result_ex_i[31:2], 2'h0 };
  assign data_addr_o_t0 = { adder_result_ex_i_t0[31:2], 2'h0 };
  assign data_we_o = lsu_we_i;
  assign data_we_o_t0 = lsu_we_i_t0;
endmodule

module auxy_noerr_rv_core_ibex(clk_i, rst_ni, clk_esc_i, rst_esc_ni, test_en_i, ram_cfg_i, hart_id_i, boot_addr_i, tl_i_o, tl_i_i, tl_d_o, tl_d_i, irq_software_i, irq_timer_i, irq_external_i, esc_tx_i, esc_rx_o, debug_req_i, crash_dump_o, lc_cpu_en_i, core_sleep_o
, tl_d_i_t0, tl_d_o_t0, boot_addr_i_t0, test_en_i_t0, esc_rx_o_t0, esc_tx_i_t0, debug_req_i_t0, hart_id_i_t0, irq_external_i_t0, irq_software_i_t0, irq_timer_i_t0, crash_dump_o_t0, core_sleep_o_t0, ram_cfg_i_t0, clk_esc_i_t0, lc_cpu_en_i_t0, rst_esc_ni_t0, tl_i_i_t0, tl_i_o_t0);
  wire [3:0] _00_;
  wire _01_;
  wire [3:0] _02_;
  wire [3:0] _03_;
  wire _04_;
  wire _05_;
  wire _06_;
  wire alert_major;
  wire alert_major_t0;
  wire alert_minor;
  wire alert_minor_t0;
  input [31:0] boot_addr_i;
  wire [31:0] boot_addr_i;
  input [31:0] boot_addr_i_t0;
  wire [31:0] boot_addr_i_t0;
  input clk_esc_i;
  wire clk_esc_i;
  input clk_esc_i_t0;
  wire clk_esc_i_t0;
  input clk_i;
  wire clk_i;
  output core_sleep_o;
  wire core_sleep_o;
  output core_sleep_o_t0;
  wire core_sleep_o_t0;
  output [127:0] crash_dump_o;
  wire [127:0] crash_dump_o;
  output [127:0] crash_dump_o_t0;
  wire [127:0] crash_dump_o_t0;
  wire [31:0] data_addr;
  wire [31:0] data_addr_t0;
  wire [3:0] data_be;
  wire [3:0] data_be_t0;
  wire data_gnt;
  wire data_gnt_t0;
  wire [31:0] data_rdata;
  wire [31:0] data_rdata_t0;
  wire data_req;
  wire data_req_t0;
  wire data_rvalid;
  wire data_rvalid_t0;
  wire [31:0] data_wdata;
  wire [31:0] data_wdata_t0;
  wire data_we;
  wire data_we_t0;
  input debug_req_i;
  wire debug_req_i;
  input debug_req_i_t0;
  wire debug_req_i_t0;
  wire esc_irq_nm;
  wire esc_irq_nm_t0;
  output [1:0] esc_rx_o;
  wire [1:0] esc_rx_o;
  output [1:0] esc_rx_o_t0;
  wire [1:0] esc_rx_o_t0;
  input [1:0] esc_tx_i;
  wire [1:0] esc_tx_i;
  input [1:0] esc_tx_i_t0;
  wire [1:0] esc_tx_i_t0;
  input [31:0] hart_id_i;
  wire [31:0] hart_id_i;
  input [31:0] hart_id_i_t0;
  wire [31:0] hart_id_i_t0;
  wire [31:0] instr_addr;
  wire [31:0] instr_addr_t0;
  wire instr_gnt;
  wire instr_gnt_t0;
  wire [31:0] instr_rdata;
  wire [31:0] instr_rdata_t0;
  wire instr_req;
  wire instr_req_t0;
  wire instr_rvalid;
  wire instr_rvalid_t0;
  input irq_external_i;
  wire irq_external_i;
  input irq_external_i_t0;
  wire irq_external_i_t0;
  wire irq_nm;
  wire irq_nm_t0;
  input irq_software_i;
  wire irq_software_i;
  input irq_software_i_t0;
  wire irq_software_i_t0;
  input irq_timer_i;
  wire irq_timer_i;
  input irq_timer_i_t0;
  wire irq_timer_i_t0;
  wire [3:0] lc_cpu_en;
  input [3:0] lc_cpu_en_i;
  wire [3:0] lc_cpu_en_i;
  input [3:0] lc_cpu_en_i_t0;
  wire [3:0] lc_cpu_en_i_t0;
  wire [3:0] lc_cpu_en_t0;
  input [9:0] ram_cfg_i;
  wire [9:0] ram_cfg_i;
  input [9:0] ram_cfg_i_t0;
  wire [9:0] ram_cfg_i_t0;
  input rst_esc_ni;
  wire rst_esc_ni;
  input rst_esc_ni_t0;
  wire rst_esc_ni_t0;
  input rst_ni;
  wire rst_ni;
  input test_en_i;
  wire test_en_i;
  input test_en_i_t0;
  wire test_en_i_t0;
  wire [65:0] tl_d_fifo2ibex;
  wire [65:0] tl_d_fifo2ibex_t0;
  input [65:0] tl_d_i;
  wire [65:0] tl_d_i;
  input [65:0] tl_d_i_t0;
  wire [65:0] tl_d_i_t0;
  wire [106:0] tl_d_ibex2fifo;
  wire [106:0] tl_d_ibex2fifo_t0;
  output [106:0] tl_d_o;
  wire [106:0] tl_d_o;
  output [106:0] tl_d_o_t0;
  wire [106:0] tl_d_o_t0;
  wire [65:0] tl_i_fifo2ibex;
  wire [65:0] tl_i_fifo2ibex_t0;
  input [65:0] tl_i_i;
  wire [65:0] tl_i_i;
  input [65:0] tl_i_i_t0;
  wire [65:0] tl_i_i_t0;
  wire [106:0] tl_i_ibex2fifo;
  wire [106:0] tl_i_ibex2fifo_t0;
  output [106:0] tl_i_o;
  wire [106:0] tl_i_o;
  output [106:0] tl_i_o_t0;
  wire [106:0] tl_i_o_t0;
  assign _01_ = | lc_cpu_en_t0;
  assign _00_ = ~ lc_cpu_en_t0;
  assign _02_ = lc_cpu_en & _00_;
  assign _03_ = 4'ha & _00_;
  assign _04_ = _02_ == _03_;
  assign _06_ = _04_ & _01_;
  assign _05_ = lc_cpu_en == 4'ha;
  paramodb54d077777a5e0334d1158f40d3ef149c7b94eb9auxy_tlul_fifo_sync  fifo_d (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .spare_req_i(1'h0),
    .spare_req_i_t0(1'h0),
    .spare_rsp_i(1'h0),
    .spare_rsp_i_t0(1'h0),
    .tl_d_i(tl_d_i),
    .tl_d_i_t0(tl_d_i_t0),
    .tl_d_o(tl_d_o),
    .tl_d_o_t0(tl_d_o_t0),
    .tl_h_i(tl_d_ibex2fifo),
    .tl_h_i_t0(tl_d_ibex2fifo_t0),
    .tl_h_o(tl_d_fifo2ibex),
    .tl_h_o_t0(tl_d_fifo2ibex_t0)
  );
  paramodb54d077777a5e0334d1158f40d3ef149c7b94eb9auxy_tlul_fifo_sync  fifo_i (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .spare_req_i(1'h0),
    .spare_req_i_t0(1'h0),
    .spare_rsp_i(1'h0),
    .spare_rsp_i_t0(1'h0),
    .tl_d_i(tl_i_i),
    .tl_d_i_t0(tl_i_i_t0),
    .tl_d_o(tl_i_o),
    .tl_d_o_t0(tl_i_o_t0),
    .tl_h_i(tl_i_ibex2fifo),
    .tl_h_i_t0(tl_i_ibex2fifo_t0),
    .tl_h_o(tl_i_fifo2ibex),
    .tl_h_o_t0(tl_i_fifo2ibex_t0)
  );
  paramodauxy_tlul_adapter_hostMAX_REQSs3200000000000000000000000000000010  tl_adapter_host_d_ibex (
    .addr_i(data_addr),
    .addr_i_t0(data_addr_t0),
    .be_i(data_be),
    .be_i_t0(data_be_t0),
    .clk_i(clk_i),
    .gnt_o(data_gnt),
    .gnt_o_t0(data_gnt_t0),
    .rdata_o(data_rdata),
    .rdata_o_t0(data_rdata_t0),
    .req_i(data_req),
    .req_i_t0(data_req_t0),
    .rst_ni(rst_ni),
    .tl_i(tl_d_fifo2ibex),
    .tl_i_t0(tl_d_fifo2ibex_t0),
    .tl_o(tl_d_ibex2fifo),
    .tl_o_t0(tl_d_ibex2fifo_t0),
    .type_i(2'h2),
    .type_i_t0(2'h0),
    .valid_o(data_rvalid),
    .valid_o_t0(data_rvalid_t0),
    .wdata_i(data_wdata),
    .wdata_i_t0(data_wdata_t0),
    .we_i(data_we),
    .we_i_t0(data_we_t0)
  );
  paramodauxy_tlul_adapter_hostMAX_REQSs3200000000000000000000000000000010  tl_adapter_host_i_ibex (
    .addr_i(instr_addr),
    .addr_i_t0(instr_addr_t0),
    .be_i(4'hf),
    .be_i_t0(4'h0),
    .clk_i(clk_i),
    .gnt_o(instr_gnt),
    .gnt_o_t0(instr_gnt_t0),
    .rdata_o(instr_rdata),
    .rdata_o_t0(instr_rdata_t0),
    .req_i(instr_req),
    .req_i_t0(instr_req_t0),
    .rst_ni(rst_ni),
    .tl_i(tl_i_fifo2ibex),
    .tl_i_t0(tl_i_fifo2ibex_t0),
    .tl_o(tl_i_ibex2fifo),
    .tl_o_t0(tl_i_ibex2fifo_t0),
    .type_i(2'h1),
    .type_i_t0(2'h0),
    .valid_o(instr_rvalid),
    .valid_o_t0(instr_rvalid_t0),
    .wdata_i(32'd0),
    .wdata_i_t0(32'd0),
    .we_i(1'h0),
    .we_i_t0(1'h0)
  );
  paramodc573af43932b4a7bfd8b52400e7bf5041b1b0ddcauxy_ibex_top  u_core (
    .alert_major_o(alert_major),
    .alert_major_o_t0(alert_major_t0),
    .alert_minor_o(alert_minor),
    .alert_minor_o_t0(alert_minor_t0),
    .boot_addr_i(boot_addr_i),
    .boot_addr_i_t0(boot_addr_i_t0),
    .clk_i(clk_i),
    .core_sleep_o(core_sleep_o),
    .core_sleep_o_t0(core_sleep_o_t0),
    .crash_dump_o(crash_dump_o),
    .crash_dump_o_t0(crash_dump_o_t0),
    .data_addr_o(data_addr),
    .data_addr_o_t0(data_addr_t0),
    .data_be_o(data_be),
    .data_be_o_t0(data_be_t0),
    .data_err_i(1'h0),
    .data_err_i_t0(1'h0),
    .data_gnt_i(data_gnt),
    .data_gnt_i_t0(data_gnt_t0),
    .data_rdata_i(data_rdata),
    .data_rdata_i_t0(data_rdata_t0),
    .data_req_o(data_req),
    .data_req_o_t0(data_req_t0),
    .data_rvalid_i(data_rvalid),
    .data_rvalid_i_t0(data_rvalid_t0),
    .data_wdata_o(data_wdata),
    .data_wdata_o_t0(data_wdata_t0),
    .data_we_o(data_we),
    .data_we_o_t0(data_we_t0),
    .debug_req_i(debug_req_i),
    .debug_req_i_t0(debug_req_i_t0),
    .fetch_enable_i(_05_),
    .fetch_enable_i_t0(_06_),
    .hart_id_i(hart_id_i),
    .hart_id_i_t0(hart_id_i_t0),
    .instr_addr_o(instr_addr),
    .instr_addr_o_t0(instr_addr_t0),
    .instr_err_i(1'h0),
    .instr_err_i_t0(1'h0),
    .instr_gnt_i(instr_gnt),
    .instr_gnt_i_t0(instr_gnt_t0),
    .instr_rdata_i(instr_rdata),
    .instr_rdata_i_t0(instr_rdata_t0),
    .instr_req_o(instr_req),
    .instr_req_o_t0(instr_req_t0),
    .instr_rvalid_i(instr_rvalid),
    .instr_rvalid_i_t0(instr_rvalid_t0),
    .irq_external_i(irq_external_i),
    .irq_external_i_t0(irq_external_i_t0),
    .irq_fast_i(15'h0000),
    .irq_fast_i_t0(15'h0000),
    .irq_nm_i(irq_nm),
    .irq_nm_i_t0(irq_nm_t0),
    .irq_software_i(irq_software_i),
    .irq_software_i_t0(irq_software_i_t0),
    .irq_timer_i(irq_timer_i),
    .irq_timer_i_t0(irq_timer_i_t0),
    .ram_cfg_i(ram_cfg_i),
    .ram_cfg_i_t0(ram_cfg_i_t0),
    .rst_ni(rst_ni),
    .test_en_i(test_en_i),
    .test_en_i_t0(test_en_i_t0)
  );
  auxy_prim_lc_sync u_lc_sync (
    .clk_i(clk_i),
    .lc_en_i(lc_cpu_en_i),
    .lc_en_i_t0(lc_cpu_en_i_t0),
    .lc_en_o(lc_cpu_en),
    .lc_en_o_t0(lc_cpu_en_t0),
    .rst_ni(rst_ni)
  );
  auxy_prim_esc_receiver u_prim_esc_receiver (
    .clk_i(clk_esc_i),
    .esc_en_o(esc_irq_nm),
    .esc_en_o_t0(esc_irq_nm_t0),
    .esc_rx_o(esc_rx_o),
    .esc_rx_o_t0(esc_rx_o_t0),
    .esc_tx_i(esc_tx_i),
    .esc_tx_i_t0(esc_tx_i_t0),
    .rst_ni(rst_esc_ni)
  );
  paramodauxy_prim_flop_2syncWidths3200000000000000000000000000000001  u_prim_flop_2sync (
    .clk_i(clk_i),
    .d_i(esc_irq_nm),
    .d_i_t0(esc_irq_nm_t0),
    .q_o(irq_nm),
    .q_o_t0(irq_nm_t0),
    .rst_ni(rst_ni)
  );
endmodule

module auxy_prim_buf(in_i, out_o, in_i_t0, out_o_t0);
  input in_i;
  wire in_i;
  input in_i_t0;
  wire in_i_t0;
  output out_o;
  wire out_o;
  output out_o_t0;
  wire out_o_t0;
  paramodauxy_prim_generic_bufWidths3200000000000000000000000000000001  \gen_generic.u_impl_generic  (
    .in_i(in_i),
    .in_i_t0(in_i_t0),
    .out_o(out_o),
    .out_o_t0(out_o_t0)
  );
endmodule

module auxy_prim_clock_gating(clk_i, en_i, test_en_i, clk_o, test_en_i_t0, en_i_t0, clk_o_t0);
  wire _00_;
  wire _01_;
  wire _02_;
  wire _03_;
  wire _04_;
  wire _05_;
  wire _06_;
  wire _07_;
  input clk_i;
  wire clk_i;
  output clk_o;
  wire clk_o;
  output clk_o_t0;
  wire clk_o_t0;
  input en_i;
  wire en_i;
  input en_i_t0;
  wire en_i_t0;
  reg en_latch;
  reg en_latch_t0;
  input test_en_i;
  wire test_en_i;
  input test_en_i_t0;
  wire test_en_i_t0;
  assign clk_o = en_latch & clk_i;
  assign clk_o_t0 = en_latch_t0 & clk_i;
  always_latch
    if (!clk_i) en_latch_t0 = _01_;
  assign _02_ = ~ en_i;
  assign _03_ = ~ test_en_i;
  assign _04_ = en_i_t0 & _03_;
  assign _05_ = test_en_i_t0 & _02_;
  assign _06_ = en_i_t0 & test_en_i_t0;
  assign _07_ = _04_ | _05_;
  assign _01_ = _07_ | _06_;
  always_latch
    if (!clk_i) en_latch = _00_;
  assign _00_ = en_i | test_en_i;
endmodule

module auxy_prim_esc_receiver(clk_i, rst_ni, esc_en_o, esc_rx_o, esc_tx_i, esc_en_o_t0, esc_rx_o_t0, esc_tx_i_t0);
  wire _000_;
  wire _001_;
  wire _002_;
  wire _003_;
  wire [2:0] _004_;
  wire [2:0] _005_;
  wire _006_;
  wire _007_;
  wire [2:0] _008_;
  wire [2:0] _009_;
  wire _010_;
  wire _011_;
  wire _012_;
  wire [2:0] _013_;
  wire [2:0] _014_;
  wire _015_;
  wire _016_;
  wire _017_;
  wire _018_;
  wire [2:0] _019_;
  wire [2:0] _020_;
  wire [2:0] _021_;
  wire [2:0] _022_;
  wire _023_;
  wire _024_;
  wire _025_;
  wire _026_;
  wire _027_;
  wire _028_;
  wire _029_;
  wire [2:0] _030_;
  wire [1:0] _031_;
  wire [2:0] _032_;
  wire _033_;
  wire _034_;
  wire _035_;
  wire _036_;
  wire _037_;
  wire [2:0] _038_;
  wire [2:0] _039_;
  wire [2:0] _040_;
  wire [2:0] _041_;
  wire [2:0] _042_;
  wire _043_;
  wire [2:0] _044_;
  wire [2:0] _045_;
  wire [2:0] _046_;
  wire _047_;
  wire _048_;
  wire _049_;
  wire _050_;
  wire _051_;
  wire _052_;
  wire _053_;
  wire _054_;
  wire _055_;
  wire [2:0] _056_;
  wire [2:0] _057_;
  wire [2:0] _058_;
  wire [2:0] _059_;
  wire [2:0] _060_;
  wire [1:0] _061_;
  wire [2:0] _062_;
  wire _063_;
  wire _064_;
  wire _065_;
  wire _066_;
  wire _067_;
  wire _068_;
  wire _069_;
  wire _070_;
  wire _071_;
  wire _072_;
  wire _073_;
  wire _074_;
  wire _075_;
  wire _076_;
  wire _077_;
  wire _078_;
  wire _079_;
  wire _080_;
  wire _081_;
  wire _082_;
  wire _083_;
  wire _084_;
  wire _085_;
  wire _086_;
  wire [2:0] _087_;
  wire [2:0] _088_;
  wire [2:0] _089_;
  wire [2:0] _090_;
  wire [2:0] _091_;
  wire [2:0] _092_;
  wire [2:0] _093_;
  wire [2:0] _094_;
  wire [2:0] _095_;
  wire [2:0] _096_;
  wire [2:0] _097_;
  wire [2:0] _098_;
  wire _099_;
  wire _100_;
  wire _101_;
  wire [2:0] _102_;
  wire [2:0] _103_;
  wire _104_;
  wire _105_;
  wire _106_;
  wire _107_;
  wire [2:0] _108_;
  wire [2:0] _109_;
  wire [2:0] _110_;
  wire _111_;
  wire _112_;
  wire _113_;
  wire [2:0] _114_;
  wire [2:0] _115_;
  wire [2:0] _116_;
  wire _117_;
  wire _118_;
  wire [2:0] _119_;
  wire [2:0] _120_;
  wire [2:0] _121_;
  wire [2:0] _122_;
  wire [2:0] _123_;
  wire _124_;
  wire _125_;
  wire [2:0] _126_;
  wire [2:0] _127_;
  wire [2:0] _128_;
  wire _129_;
  wire _130_;
  wire _131_;
  wire _132_;
  wire [2:0] _133_;
  wire [2:0] _134_;
  wire [2:0] _135_;
  wire [2:0] _136_;
  wire [2:0] _137_;
  wire _138_;
  wire _139_;
  wire _140_;
  wire _141_;
  wire _142_;
  wire _143_;
  wire _144_;
  wire _145_;
  wire _146_;
  wire _147_;
  wire _148_;
  wire _149_;
  wire [2:0] _150_;
  wire [2:0] _151_;
  wire [2:0] _152_;
  wire [2:0] _153_;
  wire [2:0] _154_;
  wire [2:0] _155_;
  wire [2:0] _156_;
  wire [2:0] _157_;
  wire [2:0] _158_;
  wire [2:0] _159_;
  wire [2:0] _160_;
  wire [2:0] _161_;
  wire _162_;
  wire _163_;
  wire [2:0] _164_;
  wire [2:0] _165_;
  wire [2:0] _166_;
  wire _167_;
  wire [2:0] _168_;
  wire [2:0] _169_;
  wire [2:0] _170_;
  wire _171_;
  wire [2:0] _172_;
  wire [2:0] _173_;
  wire [2:0] _174_;
  wire _175_;
  wire [2:0] _176_;
  wire _177_;
  wire _178_;
  wire _179_;
  wire _180_;
  wire _181_;
  wire [2:0] _182_;
  wire [2:0] _183_;
  wire [2:0] _184_;
  wire [2:0] _185_;
  wire _186_;
  wire _187_;
  wire _188_;
  wire _189_;
  wire _190_;
  wire _191_;
  wire _192_;
  wire _193_;
  wire _194_;
  wire _195_;
  wire _196_;
  wire _197_;
  wire _198_;
  wire _199_;
  wire _200_;
  wire _201_;
  wire [2:0] _202_;
  wire [2:0] _203_;
  wire [2:0] _204_;
  wire [2:0] _205_;
  wire [2:0] _206_;
  wire [2:0] _207_;
  wire _208_;
  wire _209_;
  wire _210_;
  wire _211_;
  wire _212_;
  wire _213_;
  wire _214_;
  wire _215_;
  wire _216_;
  wire _217_;
  wire _218_;
  input clk_i;
  wire clk_i;
  output esc_en_o;
  wire esc_en_o;
  output esc_en_o_t0;
  wire esc_en_o_t0;
  wire esc_level;
  wire esc_level_t0;
  output [1:0] esc_rx_o;
  wire [1:0] esc_rx_o;
  output [1:0] esc_rx_o_t0;
  wire [1:0] esc_rx_o_t0;
  input [1:0] esc_tx_i;
  wire [1:0] esc_tx_i;
  input [1:0] esc_tx_i_t0;
  wire [1:0] esc_tx_i_t0;
  wire resp_n;
  wire resp_n_t0;
  wire resp_nd;
  wire resp_nd_t0;
  reg resp_nq;
  reg resp_nq_t0;
  wire resp_p;
  wire resp_p_t0;
  wire resp_pd;
  wire resp_pd_t0;
  reg resp_pq;
  reg resp_pq_t0;
  input rst_ni;
  wire rst_ni;
  wire sigint_detected;
  wire sigint_detected_t0;
  wire [2:0] state_d;
  wire [2:0] state_d_t0;
  reg [2:0] state_q;
  reg [2:0] state_q_t0;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) resp_pq_t0 <= 1'h0;
    else resp_pq_t0 <= resp_pd_t0;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) resp_nq_t0 <= 1'h0;
    else resp_nq_t0 <= resp_nd_t0;
  assign _029_ = ~ _023_;
  assign _176_ = state_d ^ state_q;
  assign _133_ = state_d_t0 | state_q_t0;
  assign _134_ = _176_ | _133_;
  assign _056_ = { _023_, _023_, _023_ } & state_d_t0;
  assign _057_ = { _029_, _029_, _029_ } & state_q_t0;
  assign _058_ = _134_ & { _024_, _024_, _024_ };
  assign _135_ = _056_ | _057_;
  assign _136_ = _135_ | _058_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) state_q_t0 <= 3'h0;
    else state_q_t0 <= _136_;
  assign _049_ = | { _137_[2:1], esc_level_t0 };
  assign _052_ = | state_q_t0;
  assign _030_ = ~ { _137_[2:1], esc_level_t0 };
  assign _042_ = ~ state_q_t0;
  assign _059_ = { _218_, _208_, esc_level } & _030_;
  assign _102_ = state_q & _042_;
  assign _060_ = 3'h4 & _030_;
  assign _103_ = 3'h4 & _042_;
  assign _126_ = 3'h3 & _042_;
  assign _127_ = 3'h2 & _042_;
  assign _128_ = 3'h1 & _042_;
  assign _186_ = _059_ == _060_;
  assign _187_ = _102_ == _103_;
  assign _188_ = _102_ == _126_;
  assign _189_ = _102_ == _127_;
  assign _190_ = _102_ == _128_;
  assign _024_ = _186_ & _049_;
  assign _210_ = _187_ & _052_;
  assign _213_ = _188_ & _052_;
  assign _215_ = _189_ & _052_;
  assign _217_ = _190_ & _052_;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) state_q <= 3'h0;
    else if (_023_) state_q <= state_d;
  assign _099_ = sigint_detected_t0 & _209_;
  assign _100_ = _210_ & sigint_detected;
  assign _101_ = sigint_detected_t0 & _210_;
  assign _162_ = _099_ | _100_;
  assign _137_[1] = _162_ | _101_;
  assign _050_ = | { _215_, _213_ };
  assign _051_ = | { _217_, _215_, _213_ };
  assign _031_ = ~ { _215_, _213_ };
  assign _032_ = ~ { _217_, _215_, _213_ };
  assign _061_ = { _214_, _212_ } & _031_;
  assign _062_ = { _216_, _214_, _212_ } & _032_;
  assign _053_ = ! _061_;
  assign _054_ = ! _062_;
  assign _055_ = ! _102_;
  assign _026_ = _053_ & _050_;
  assign _028_ = _054_ & _051_;
  assign _137_[2] = _055_ & _052_;
  assign _034_ = ~ _211_;
  assign _036_ = ~ _214_;
  assign _037_ = ~ _129_;
  assign _038_ = ~ { _211_, _211_, _211_ };
  assign _039_ = ~ { _218_, _218_, _218_ };
  assign _040_ = ~ { _216_, _216_, _216_ };
  assign _041_ = ~ { _131_, _131_, _131_ };
  assign _043_ = ~ _208_;
  assign _044_ = ~ { _208_, _208_, _208_ };
  assign _045_ = ~ { sigint_detected, sigint_detected, sigint_detected };
  assign _046_ = ~ { esc_level, esc_level, esc_level };
  assign _140_ = _210_ | _034_;
  assign _144_ = _215_ | _036_;
  assign _145_ = _130_ | _037_;
  assign _150_ = { _210_, _210_, _210_ } | _038_;
  assign _153_ = { _137_[2], _137_[2], _137_[2] } | _039_;
  assign _156_ = { _217_, _217_, _217_ } | _040_;
  assign _159_ = { _132_, _132_, _132_ } | _041_;
  assign _163_ = _137_[1] | _043_;
  assign _164_ = { _137_[1], _137_[1], _137_[1] } | _044_;
  assign _168_ = { sigint_detected_t0, sigint_detected_t0, sigint_detected_t0 } | _045_;
  assign _172_ = { esc_level_t0, esc_level_t0, esc_level_t0 } | _046_;
  assign _141_ = _210_ | _211_;
  assign _143_ = _137_[2] | _218_;
  assign _146_ = _130_ | _129_;
  assign _151_ = { _210_, _210_, _210_ } | { _211_, _211_, _211_ };
  assign _154_ = { _137_[2], _137_[2], _137_[2] } | { _218_, _218_, _218_ };
  assign _157_ = { _217_, _217_, _217_ } | { _216_, _216_, _216_ };
  assign _160_ = { _132_, _132_, _132_ } | { _131_, _131_, _131_ };
  assign _165_ = { _137_[1], _137_[1], _137_[1] } | { _208_, _208_, _208_ };
  assign _167_ = sigint_detected_t0 | sigint_detected;
  assign _169_ = { sigint_detected_t0, sigint_detected_t0, sigint_detected_t0 } | { sigint_detected, sigint_detected, sigint_detected };
  assign _171_ = esc_level_t0 | esc_level;
  assign _173_ = { esc_level_t0, esc_level_t0, esc_level_t0 } | { esc_level, esc_level, esc_level };
  assign _175_ = _028_ | _027_;
  assign _074_ = _193_ & _144_;
  assign _076_ = _195_ & _145_;
  assign _069_ = _011_ & _140_;
  assign _082_ = _199_ & _144_;
  assign _084_ = _201_ & _145_;
  assign _087_ = _020_ & _150_;
  assign _090_ = 3'h0 & _153_;
  assign _093_ = _205_ & _156_;
  assign _096_ = _207_ & _159_;
  assign _104_ = _001_ & _163_;
  assign _106_ = _003_ & _163_;
  assign _108_ = _005_ & _164_;
  assign _114_ = 3'h0 & _168_;
  assign _119_ = 3'h0 & _172_;
  assign _070_ = _016_ & _141_;
  assign _077_ = _192_ & _146_;
  assign _079_ = _018_ & _141_;
  assign _072_ = esc_level_t0 & _143_;
  assign _085_ = _197_ & _146_;
  assign _088_ = _022_ & _151_;
  assign _091_ = _009_ & _154_;
  assign _094_ = _014_ & _157_;
  assign _097_ = _203_ & _160_;
  assign _109_ = 3'h0 & _165_;
  assign _111_ = resp_pq_t0 & _167_;
  assign _115_ = 3'h0 & _169_;
  assign _117_ = resp_pq_t0 & _171_;
  assign _120_ = 3'h0 & _173_;
  assign _124_ = esc_level_t0 & _175_;
  assign _142_ = _069_ | _070_;
  assign _147_ = _076_ | _077_;
  assign _148_ = _069_ | _079_;
  assign _149_ = _084_ | _085_;
  assign _152_ = _087_ | _088_;
  assign _155_ = _090_ | _091_;
  assign _158_ = _093_ | _094_;
  assign _161_ = _096_ | _097_;
  assign _166_ = _108_ | _109_;
  assign _170_ = _114_ | _115_;
  assign _174_ = _119_ | _120_;
  assign _177_ = _010_ ^ _015_;
  assign _179_ = _194_ ^ _191_;
  assign _180_ = _012_ ^ _017_;
  assign _181_ = _200_ ^ _196_;
  assign _182_ = _019_ ^ _021_;
  assign _183_ = _204_ ^ _013_;
  assign _184_ = _206_ ^ _202_;
  assign _185_ = _004_ ^ 3'h4;
  assign _071_ = _210_ & _177_;
  assign _073_ = _137_[2] & esc_level;
  assign _075_ = _215_ & _178_;
  assign _078_ = _130_ & _179_;
  assign _080_ = _210_ & _180_;
  assign _081_ = _137_[2] & _006_;
  assign _083_ = _215_ & _047_;
  assign _086_ = _130_ & _181_;
  assign _089_ = { _210_, _210_, _210_ } & _182_;
  assign _092_ = { _137_[2], _137_[2], _137_[2] } & _008_;
  assign _095_ = { _217_, _217_, _217_ } & _183_;
  assign _098_ = { _132_, _132_, _132_ } & _184_;
  assign _105_ = _137_[1] & _000_;
  assign _107_ = _137_[1] & _002_;
  assign _110_ = { _137_[1], _137_[1], _137_[1] } & _185_;
  assign _112_ = sigint_detected_t0 & resp_pq;
  assign _113_ = sigint_detected_t0 & _048_;
  assign _116_ = { sigint_detected_t0, sigint_detected_t0, sigint_detected_t0 } & 3'h4;
  assign _118_ = esc_level_t0 & _048_;
  assign _121_ = { esc_level_t0, esc_level_t0, esc_level_t0 } & 3'h3;
  assign _122_ = { esc_level_t0, esc_level_t0, esc_level_t0 } & 3'h1;
  assign _123_ = { esc_level_t0, esc_level_t0, esc_level_t0 } & 3'hx;
  assign _125_ = _028_ & _006_;
  assign _192_ = _071_ | _142_;
  assign _193_ = _073_ | _072_;
  assign _195_ = _075_ | _074_;
  assign _001_ = _078_ | _147_;
  assign _197_ = _080_ | _148_;
  assign _199_ = _081_ | _072_;
  assign _201_ = _083_ | _082_;
  assign _003_ = _086_ | _149_;
  assign _203_ = _089_ | _152_;
  assign _205_ = _092_ | _155_;
  assign _207_ = _095_ | _158_;
  assign _005_ = _098_ | _161_;
  assign resp_n_t0 = _105_ | _104_;
  assign resp_p_t0 = _107_ | _106_;
  assign state_d_t0 = _110_ | _166_;
  assign _016_ = _112_ | _111_;
  assign _018_ = _113_ | _111_;
  assign _022_ = _116_ | _170_;
  assign _011_ = _118_ | _117_;
  assign _020_ = _121_ | _174_;
  assign _014_ = _122_ | _174_;
  assign _009_ = _123_ | _174_;
  assign esc_en_o_t0 = _125_ | _124_;
  assign _023_ = { _218_, _208_, esc_level } != 3'h4;
  assign _047_ = ~ _198_;
  assign _048_ = ~ resp_pq;
  assign _025_ = | { _214_, _212_ };
  assign _027_ = | { _216_, _214_, _212_ };
  assign _033_ = ~ _212_;
  assign _035_ = ~ _025_;
  assign _063_ = _213_ & _034_;
  assign _066_ = _026_ & _034_;
  assign _064_ = _210_ & _033_;
  assign _067_ = _210_ & _035_;
  assign _065_ = _213_ & _210_;
  assign _068_ = _026_ & _210_;
  assign _138_ = _063_ | _064_;
  assign _139_ = _066_ | _067_;
  assign _130_ = _138_ | _065_;
  assign _132_ = _139_ | _068_;
  assign _129_ = _212_ | _211_;
  assign _131_ = _025_ | _211_;
  assign _191_ = _211_ ? _015_ : _010_;
  assign _178_ = _218_ ? _007_ : 1'h1;
  assign _194_ = _214_ ? 1'h0 : _178_;
  assign _000_ = _129_ ? _191_ : _194_;
  assign _196_ = _211_ ? _017_ : _012_;
  assign _198_ = _218_ ? _006_ : 1'h0;
  assign _200_ = _214_ ? 1'h1 : _198_;
  assign _002_ = _129_ ? _196_ : _200_;
  assign _202_ = _211_ ? _021_ : _019_;
  assign _204_ = _218_ ? _008_ : 3'h0;
  assign _206_ = _216_ ? _013_ : _204_;
  assign _004_ = _131_ ? _202_ : _206_;
  assign _208_ = sigint_detected && _209_;
  assign _209_ = state_q != 3'h4;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) resp_pq <= 1'h0;
    else resp_pq <= resp_pd;
  always_ff @(posedge clk_i, negedge rst_ni)
    if (!rst_ni) resp_nq <= 1'h1;
    else resp_nq <= resp_nd;
  assign resp_n = _208_ ? 1'h0 : _000_;
  assign resp_p = _208_ ? 1'h0 : _002_;
  assign state_d = _208_ ? 3'h4 : _004_;
  assign _015_ = sigint_detected ? _048_ : 1'h1;
  assign _017_ = sigint_detected ? _048_ : 1'h0;
  assign _021_ = sigint_detected ? 3'h4 : 3'h0;
  assign _010_ = esc_level ? resp_pq : 1'h1;
  assign _012_ = esc_level ? _048_ : 1'h0;
  assign _019_ = esc_level ? 3'h3 : 3'h0;
  assign _006_ = esc_level ? 1'h1 : 1'h0;
  assign _013_ = esc_level ? 3'h3 : 3'h2;
  assign _007_ = esc_level ? 1'h0 : 1'h1;
  assign _008_ = esc_level ? 3'h1 : 3'hx;
  assign _211_ = state_q == 3'h4;
  assign _218_ = ! state_q;
  assign esc_en_o = _027_ ? _006_ : 1'h0;
  assign _212_ = state_q == 3'h3;
  assign _214_ = state_q == 3'h2;
  assign _216_ = state_q == 3'h1;
  paramodauxy_prim_diff_decodeAsyncOn10  i_decode_esc (
    .clk_i(clk_i),
    .diff_ni(esc_tx_i[0]),
    .diff_ni_t0(esc_tx_i_t0[0]),
    .diff_pi(esc_tx_i[1]),
    .diff_pi_t0(esc_tx_i_t0[1]),
    .level_o(esc_level),
    .level_o_t0(esc_level_t0),
    .rst_ni(rst_ni),
    .sigint_o(sigint_detected),
    .sigint_o_t0(sigint_detected_t0)
  );
  auxy_prim_buf u_prim_buf_n (
    .in_i(resp_n),
    .in_i_t0(resp_n_t0),
    .out_o(resp_nd),
    .out_o_t0(resp_nd_t0)
  );
  auxy_prim_buf u_prim_buf_p (
    .in_i(resp_p),
    .in_i_t0(resp_p_t0),
    .out_o(resp_pd),
    .out_o_t0(resp_pd_t0)
  );
  assign _137_[0] = esc_level_t0;
  assign esc_rx_o = { resp_pq, resp_nq };
  assign esc_rx_o_t0 = { resp_pq_t0, resp_nq_t0 };
endmodule

module auxy_prim_lc_sync(clk_i, rst_ni, lc_en_i, lc_en_o, lc_en_o_t0, lc_en_i_t0);
  input clk_i;
  wire clk_i;
  wire [3:0] lc_en;
  input [3:0] lc_en_i;
  wire [3:0] lc_en_i;
  input [3:0] lc_en_i_t0;
  wire [3:0] lc_en_i_t0;
  output [3:0] lc_en_o;
  wire [3:0] lc_en_o;
  output [3:0] lc_en_o_t0;
  wire [3:0] lc_en_o_t0;
  wire [3:0] lc_en_t0;
  input rst_ni;
  wire rst_ni;
  auxy_prim_buf \gen_buffs[0].gen_bits[0].u_prim_buf  (
    .in_i(lc_en[0]),
    .in_i_t0(lc_en_t0[0]),
    .out_o(lc_en_o[0]),
    .out_o_t0(lc_en_o_t0[0])
  );
  auxy_prim_buf \gen_buffs[0].gen_bits[1].u_prim_buf  (
    .in_i(lc_en[1]),
    .in_i_t0(lc_en_t0[1]),
    .out_o(lc_en_o[1]),
    .out_o_t0(lc_en_o_t0[1])
  );
  auxy_prim_buf \gen_buffs[0].gen_bits[2].u_prim_buf  (
    .in_i(lc_en[2]),
    .in_i_t0(lc_en_t0[2]),
    .out_o(lc_en_o[2]),
    .out_o_t0(lc_en_o_t0[2])
  );
  auxy_prim_buf \gen_buffs[0].gen_bits[3].u_prim_buf  (
    .in_i(lc_en[3]),
    .in_i_t0(lc_en_t0[3]),
    .out_o(lc_en_o[3]),
    .out_o_t0(lc_en_o_t0[3])
  );
  paramod6ae18350b51be32fd7406c5aaac3c7582e0e6af0auxy_prim_flop_2sync  \gen_flops.u_prim_flop_2sync  (
    .clk_i(clk_i),
    .d_i(lc_en_i),
    .d_i_t0(lc_en_i_t0),
    .q_o(lc_en),
    .q_o_t0(lc_en_t0),
    .rst_ni(rst_ni)
  );
endmodule

module auxy_prim_secded_64_57_dec(in, d_o, syndrome_o, err_o, err_o_t0, in_t0, d_o_t0, syndrome_o_t0);
  wire [63:0] _000_;
  wire [63:0] _001_;
  wire [63:0] _002_;
  wire [63:0] _003_;
  wire [63:0] _004_;
  wire [63:0] _005_;
  wire [63:0] _006_;
  wire [63:0] _007_;
  wire [63:0] _008_;
  wire [63:0] _009_;
  wire [63:0] _010_;
  wire [63:0] _011_;
  wire [63:0] _012_;
  wire [63:0] _013_;
  wire [6:0] _014_;
  wire _015_;
  wire [63:0] _016_;
  wire [63:0] _017_;
  wire [63:0] _018_;
  wire [63:0] _019_;
  wire [63:0] _020_;
  wire [63:0] _021_;
  wire [63:0] _022_;
  wire [63:0] _023_;
  wire [63:0] _024_;
  wire _025_;
  wire _026_;
  wire _027_;
  wire [6:0] _028_;
  wire [6:0] _029_;
  wire [6:0] _030_;
  wire [6:0] _031_;
  wire [6:0] _032_;
  wire [6:0] _033_;
  wire [6:0] _034_;
  wire [6:0] _035_;
  wire [6:0] _036_;
  wire [6:0] _037_;
  wire [6:0] _038_;
  wire [6:0] _039_;
  wire [6:0] _040_;
  wire [6:0] _041_;
  wire [6:0] _042_;
  wire [6:0] _043_;
  wire [6:0] _044_;
  wire [6:0] _045_;
  wire [6:0] _046_;
  wire [6:0] _047_;
  wire [6:0] _048_;
  wire [6:0] _049_;
  wire [6:0] _050_;
  wire [6:0] _051_;
  wire [6:0] _052_;
  wire [6:0] _053_;
  wire [6:0] _054_;
  wire [6:0] _055_;
  wire [6:0] _056_;
  wire [6:0] _057_;
  wire [6:0] _058_;
  wire [6:0] _059_;
  wire [6:0] _060_;
  wire [6:0] _061_;
  wire [6:0] _062_;
  wire [6:0] _063_;
  wire [6:0] _064_;
  wire [6:0] _065_;
  wire [6:0] _066_;
  wire [6:0] _067_;
  wire [6:0] _068_;
  wire [6:0] _069_;
  wire [6:0] _070_;
  wire [6:0] _071_;
  wire [6:0] _072_;
  wire [6:0] _073_;
  wire [6:0] _074_;
  wire [6:0] _075_;
  wire [6:0] _076_;
  wire [6:0] _077_;
  wire [6:0] _078_;
  wire [6:0] _079_;
  wire [6:0] _080_;
  wire [6:0] _081_;
  wire [6:0] _082_;
  wire [6:0] _083_;
  wire [6:0] _084_;
  wire [6:0] _085_;
  wire [63:0] _086_;
  wire [63:0] _087_;
  wire [63:0] _088_;
  wire [63:0] _089_;
  wire [63:0] _090_;
  wire [63:0] _091_;
  wire [63:0] _092_;
  wire _093_;
  wire _094_;
  wire _095_;
  wire _096_;
  wire _097_;
  wire _098_;
  wire _099_;
  wire _100_;
  wire _101_;
  wire _102_;
  wire _103_;
  wire _104_;
  wire _105_;
  wire _106_;
  wire _107_;
  wire _108_;
  wire _109_;
  wire _110_;
  wire _111_;
  wire _112_;
  wire _113_;
  wire _114_;
  wire _115_;
  wire _116_;
  wire _117_;
  wire _118_;
  wire _119_;
  wire _120_;
  wire _121_;
  wire _122_;
  wire _123_;
  wire _124_;
  wire _125_;
  wire _126_;
  wire _127_;
  wire _128_;
  wire _129_;
  wire _130_;
  wire _131_;
  wire _132_;
  wire _133_;
  wire _134_;
  wire _135_;
  wire _136_;
  wire _137_;
  wire _138_;
  wire _139_;
  wire _140_;
  wire _141_;
  wire _142_;
  wire _143_;
  wire _144_;
  wire _145_;
  wire _146_;
  wire _147_;
  wire _148_;
  wire _149_;
  wire _150_;
  wire _151_;
  wire _152_;
  wire _153_;
  wire _154_;
  wire _155_;
  wire _156_;
  wire _157_;
  wire _158_;
  wire _159_;
  wire _160_;
  wire _161_;
  wire _162_;
  wire _163_;
  wire _164_;
  wire _165_;
  wire _166_;
  wire _167_;
  wire _168_;
  wire _169_;
  wire _170_;
  wire _171_;
  wire _172_;
  wire _173_;
  wire _174_;
  wire _175_;
  wire _176_;
  wire _177_;
  wire _178_;
  wire _179_;
  wire _180_;
  wire _181_;
  wire _182_;
  wire _183_;
  wire _184_;
  wire _185_;
  wire _186_;
  wire _187_;
  wire _188_;
  wire _189_;
  wire _190_;
  wire _191_;
  wire _192_;
  wire _193_;
  wire _194_;
  wire _195_;
  wire _196_;
  wire _197_;
  wire _198_;
  wire _199_;
  wire _200_;
  wire _201_;
  wire _202_;
  wire _203_;
  wire _204_;
  wire _205_;
  wire _206_;
  wire _207_;
  wire _208_;
  wire _209_;
  wire _210_;
  wire _211_;
  wire _212_;
  wire _213_;
  wire _214_;
  wire _215_;
  wire _216_;
  wire _217_;
  wire _218_;
  wire _219_;
  wire _220_;
  wire _221_;
  wire _222_;
  wire _223_;
  wire _224_;
  wire _225_;
  wire _226_;
  wire _227_;
  wire _228_;
  wire _229_;
  wire _230_;
  wire _231_;
  wire _232_;
  wire _233_;
  wire _234_;
  wire _235_;
  wire _236_;
  wire _237_;
  wire _238_;
  wire _239_;
  wire _240_;
  wire _241_;
  wire _242_;
  wire _243_;
  wire _244_;
  wire _245_;
  wire _246_;
  wire _247_;
  wire _248_;
  wire _249_;
  wire _250_;
  wire _251_;
  wire _252_;
  wire _253_;
  wire _254_;
  wire _255_;
  wire _256_;
  wire _257_;
  wire _258_;
  wire _259_;
  wire _260_;
  wire _261_;
  wire _262_;
  wire _263_;
  wire _264_;
  wire _265_;
  wire _266_;
  wire _267_;
  output [56:0] d_o;
  wire [56:0] d_o;
  output [56:0] d_o_t0;
  wire [56:0] d_o_t0;
  output [1:0] err_o;
  wire [1:0] err_o;
  output [1:0] err_o_t0;
  wire [1:0] err_o_t0;
  input [63:0] in;
  wire [63:0] in;
  input [63:0] in_t0;
  wire [63:0] in_t0;
  wire single_error;
  wire single_error_t0;
  output [6:0] syndrome_o;
  wire [6:0] syndrome_o;
  output [6:0] syndrome_o_t0;
  wire [6:0] syndrome_o_t0;
  assign _000_ = in & 64'h0303fff800007fff;
  assign _002_ = in & 64'h057c1ff801ff801f;
  assign _004_ = in & 64'h09bde1f87e0781e1;
  assign _006_ = in & 64'h11deee3b8e388e22;
  assign _008_ = in & 64'h21ef76cdb2c93244;
  assign _010_ = in & 64'h41f7bb56d5525488;
  assign _012_ = in & 64'h81fbdda769a46910;
  assign err_o[1] = _265_ & _266_;
  assign _016_ = in_t0 & 64'h0303fff800007fff;
  assign _019_ = in_t0 & 64'h057c1ff801ff801f;
  assign _020_ = in_t0 & 64'h09bde1f87e0781e1;
  assign _021_ = in_t0 & 64'h11deee3b8e388e22;
  assign _022_ = in_t0 & 64'h21ef76cdb2c93244;
  assign _023_ = in_t0 & 64'h41f7bb56d5525488;
  assign _024_ = in_t0 & 64'h81fbdda769a46910;
  assign _025_ = single_error_t0 & _266_;
  assign _017_ = 64'h0000000000000000 & in;
  assign _026_ = _267_ & _265_;
  assign _018_ = in_t0 & 64'h0000000000000000;
  assign _027_ = single_error_t0 & _267_;
  assign _086_ = _016_ | _017_;
  assign _087_ = _019_ | _017_;
  assign _088_ = _020_ | _017_;
  assign _089_ = _021_ | _017_;
  assign _090_ = _022_ | _017_;
  assign _091_ = _023_ | _017_;
  assign _092_ = _024_ | _017_;
  assign _093_ = _025_ | _026_;
  assign _001_ = _086_ | _018_;
  assign _003_ = _087_ | _018_;
  assign _005_ = _088_ | _018_;
  assign _007_ = _089_ | _018_;
  assign _009_ = _090_ | _018_;
  assign _011_ = _091_ | _018_;
  assign _013_ = _092_ | _018_;
  assign err_o_t0[1] = _093_ | _027_;
  assign _014_ = ~ syndrome_o_t0;
  assign _028_ = syndrome_o & _014_;
  assign _029_ = 7'h07 & _014_;
  assign _030_ = 7'h0b & _014_;
  assign _031_ = 7'h13 & _014_;
  assign _032_ = 7'h23 & _014_;
  assign _033_ = 7'h43 & _014_;
  assign _034_ = 7'h0d & _014_;
  assign _035_ = 7'h15 & _014_;
  assign _036_ = 7'h25 & _014_;
  assign _037_ = 7'h45 & _014_;
  assign _038_ = 7'h19 & _014_;
  assign _039_ = 7'h29 & _014_;
  assign _040_ = 7'h49 & _014_;
  assign _041_ = 7'h31 & _014_;
  assign _042_ = 7'h51 & _014_;
  assign _043_ = 7'h61 & _014_;
  assign _044_ = 7'h0e & _014_;
  assign _045_ = 7'h16 & _014_;
  assign _046_ = 7'h26 & _014_;
  assign _047_ = 7'h46 & _014_;
  assign _048_ = 7'h1a & _014_;
  assign _049_ = 7'h2a & _014_;
  assign _050_ = 7'h4a & _014_;
  assign _051_ = 7'h32 & _014_;
  assign _052_ = 7'h52 & _014_;
  assign _053_ = 7'h62 & _014_;
  assign _054_ = 7'h1c & _014_;
  assign _055_ = 7'h2c & _014_;
  assign _056_ = 7'h4c & _014_;
  assign _057_ = 7'h34 & _014_;
  assign _058_ = 7'h54 & _014_;
  assign _059_ = 7'h64 & _014_;
  assign _060_ = 7'h38 & _014_;
  assign _061_ = 7'h58 & _014_;
  assign _062_ = 7'h68 & _014_;
  assign _063_ = 7'h70 & _014_;
  assign _064_ = 7'h1f & _014_;
  assign _065_ = 7'h2f & _014_;
  assign _066_ = 7'h4f & _014_;
  assign _067_ = 7'h37 & _014_;
  assign _068_ = 7'h57 & _014_;
  assign _069_ = 7'h67 & _014_;
  assign _070_ = 7'h3b & _014_;
  assign _071_ = 7'h5b & _014_;
  assign _072_ = 7'h6b & _014_;
  assign _073_ = 7'h73 & _014_;
  assign _074_ = 7'h3d & _014_;
  assign _075_ = 7'h5d & _014_;
  assign _076_ = 7'h6d & _014_;
  assign _077_ = 7'h75 & _014_;
  assign _078_ = 7'h79 & _014_;
  assign _079_ = 7'h3e & _014_;
  assign _080_ = 7'h5e & _014_;
  assign _081_ = 7'h6e & _014_;
  assign _082_ = 7'h76 & _014_;
  assign _083_ = 7'h7a & _014_;
  assign _084_ = 7'h7c & _014_;
  assign _085_ = 7'h7f & _014_;
  assign _094_ = _028_ == _029_;
  assign _095_ = _028_ == _030_;
  assign _096_ = _028_ == _031_;
  assign _097_ = _028_ == _032_;
  assign _098_ = _028_ == _033_;
  assign _099_ = _028_ == _034_;
  assign _100_ = _028_ == _035_;
  assign _101_ = _028_ == _036_;
  assign _102_ = _028_ == _037_;
  assign _103_ = _028_ == _038_;
  assign _104_ = _028_ == _039_;
  assign _105_ = _028_ == _040_;
  assign _106_ = _028_ == _041_;
  assign _107_ = _028_ == _042_;
  assign _108_ = _028_ == _043_;
  assign _109_ = _028_ == _044_;
  assign _110_ = _028_ == _045_;
  assign _111_ = _028_ == _046_;
  assign _112_ = _028_ == _047_;
  assign _113_ = _028_ == _048_;
  assign _114_ = _028_ == _049_;
  assign _115_ = _028_ == _050_;
  assign _116_ = _028_ == _051_;
  assign _117_ = _028_ == _052_;
  assign _118_ = _028_ == _053_;
  assign _119_ = _028_ == _054_;
  assign _120_ = _028_ == _055_;
  assign _121_ = _028_ == _056_;
  assign _122_ = _028_ == _057_;
  assign _123_ = _028_ == _058_;
  assign _124_ = _028_ == _059_;
  assign _125_ = _028_ == _060_;
  assign _126_ = _028_ == _061_;
  assign _127_ = _028_ == _062_;
  assign _128_ = _028_ == _063_;
  assign _129_ = _028_ == _064_;
  assign _130_ = _028_ == _065_;
  assign _131_ = _028_ == _066_;
  assign _132_ = _028_ == _067_;
  assign _133_ = _028_ == _068_;
  assign _134_ = _028_ == _069_;
  assign _135_ = _028_ == _070_;
  assign _136_ = _028_ == _071_;
  assign _137_ = _028_ == _072_;
  assign _138_ = _028_ == _073_;
  assign _139_ = _028_ == _074_;
  assign _140_ = _028_ == _075_;
  assign _141_ = _028_ == _076_;
  assign _142_ = _028_ == _077_;
  assign _143_ = _028_ == _078_;
  assign _144_ = _028_ == _079_;
  assign _145_ = _028_ == _080_;
  assign _146_ = _028_ == _081_;
  assign _147_ = _028_ == _082_;
  assign _148_ = _028_ == _083_;
  assign _149_ = _028_ == _084_;
  assign _150_ = _028_ == _085_;
  assign _152_ = _094_ & single_error_t0;
  assign _154_ = _095_ & single_error_t0;
  assign _156_ = _096_ & single_error_t0;
  assign _158_ = _097_ & single_error_t0;
  assign _160_ = _098_ & single_error_t0;
  assign _162_ = _099_ & single_error_t0;
  assign _164_ = _100_ & single_error_t0;
  assign _166_ = _101_ & single_error_t0;
  assign _168_ = _102_ & single_error_t0;
  assign _170_ = _103_ & single_error_t0;
  assign _172_ = _104_ & single_error_t0;
  assign _174_ = _105_ & single_error_t0;
  assign _176_ = _106_ & single_error_t0;
  assign _178_ = _107_ & single_error_t0;
  assign _180_ = _108_ & single_error_t0;
  assign _182_ = _109_ & single_error_t0;
  assign _184_ = _110_ & single_error_t0;
  assign _186_ = _111_ & single_error_t0;
  assign _188_ = _112_ & single_error_t0;
  assign _190_ = _113_ & single_error_t0;
  assign _192_ = _114_ & single_error_t0;
  assign _194_ = _115_ & single_error_t0;
  assign _196_ = _116_ & single_error_t0;
  assign _198_ = _117_ & single_error_t0;
  assign _200_ = _118_ & single_error_t0;
  assign _202_ = _119_ & single_error_t0;
  assign _204_ = _120_ & single_error_t0;
  assign _206_ = _121_ & single_error_t0;
  assign _208_ = _122_ & single_error_t0;
  assign _210_ = _123_ & single_error_t0;
  assign _212_ = _124_ & single_error_t0;
  assign _214_ = _125_ & single_error_t0;
  assign _216_ = _126_ & single_error_t0;
  assign _218_ = _127_ & single_error_t0;
  assign _220_ = _128_ & single_error_t0;
  assign _222_ = _129_ & single_error_t0;
  assign _224_ = _130_ & single_error_t0;
  assign _226_ = _131_ & single_error_t0;
  assign _228_ = _132_ & single_error_t0;
  assign _230_ = _133_ & single_error_t0;
  assign _232_ = _134_ & single_error_t0;
  assign _234_ = _135_ & single_error_t0;
  assign _236_ = _136_ & single_error_t0;
  assign _238_ = _137_ & single_error_t0;
  assign _240_ = _138_ & single_error_t0;
  assign _242_ = _139_ & single_error_t0;
  assign _244_ = _140_ & single_error_t0;
  assign _246_ = _141_ & single_error_t0;
  assign _248_ = _142_ & single_error_t0;
  assign _250_ = _143_ & single_error_t0;
  assign _252_ = _144_ & single_error_t0;
  assign _254_ = _145_ & single_error_t0;
  assign _256_ = _146_ & single_error_t0;
  assign _258_ = _147_ & single_error_t0;
  assign _260_ = _148_ & single_error_t0;
  assign _262_ = _149_ & single_error_t0;
  assign _264_ = _150_ & single_error_t0;
  assign _015_ = ! _028_;
  assign _267_ = _015_ & single_error_t0;
  assign syndrome_o_t0[0] = | _001_;
  assign syndrome_o_t0[1] = | _003_;
  assign syndrome_o_t0[2] = | _005_;
  assign syndrome_o_t0[3] = | _007_;
  assign syndrome_o_t0[4] = | _009_;
  assign syndrome_o_t0[5] = | _011_;
  assign syndrome_o_t0[6] = | _013_;
  assign single_error_t0 = | { _013_, _011_, _009_, _007_, _005_, _003_, _001_ };
  assign d_o_t0[0] = _152_ | in_t0[0];
  assign d_o_t0[1] = _154_ | in_t0[1];
  assign d_o_t0[2] = _156_ | in_t0[2];
  assign d_o_t0[3] = _158_ | in_t0[3];
  assign d_o_t0[4] = _160_ | in_t0[4];
  assign d_o_t0[5] = _162_ | in_t0[5];
  assign d_o_t0[6] = _164_ | in_t0[6];
  assign d_o_t0[7] = _166_ | in_t0[7];
  assign d_o_t0[8] = _168_ | in_t0[8];
  assign d_o_t0[9] = _170_ | in_t0[9];
  assign d_o_t0[10] = _172_ | in_t0[10];
  assign d_o_t0[11] = _174_ | in_t0[11];
  assign d_o_t0[12] = _176_ | in_t0[12];
  assign d_o_t0[13] = _178_ | in_t0[13];
  assign d_o_t0[14] = _180_ | in_t0[14];
  assign d_o_t0[15] = _182_ | in_t0[15];
  assign d_o_t0[16] = _184_ | in_t0[16];
  assign d_o_t0[17] = _186_ | in_t0[17];
  assign d_o_t0[18] = _188_ | in_t0[18];
  assign d_o_t0[19] = _190_ | in_t0[19];
  assign d_o_t0[20] = _192_ | in_t0[20];
  assign d_o_t0[21] = _194_ | in_t0[21];
  assign d_o_t0[22] = _196_ | in_t0[22];
  assign d_o_t0[23] = _198_ | in_t0[23];
  assign d_o_t0[24] = _200_ | in_t0[24];
  assign d_o_t0[25] = _202_ | in_t0[25];
  assign d_o_t0[26] = _204_ | in_t0[26];
  assign d_o_t0[27] = _206_ | in_t0[27];
  assign d_o_t0[28] = _208_ | in_t0[28];
  assign d_o_t0[29] = _210_ | in_t0[29];
  assign d_o_t0[30] = _212_ | in_t0[30];
  assign d_o_t0[31] = _214_ | in_t0[31];
  assign d_o_t0[32] = _216_ | in_t0[32];
  assign d_o_t0[33] = _218_ | in_t0[33];
  assign d_o_t0[34] = _220_ | in_t0[34];
  assign d_o_t0[35] = _222_ | in_t0[35];
  assign d_o_t0[36] = _224_ | in_t0[36];
  assign d_o_t0[37] = _226_ | in_t0[37];
  assign d_o_t0[38] = _228_ | in_t0[38];
  assign d_o_t0[39] = _230_ | in_t0[39];
  assign d_o_t0[40] = _232_ | in_t0[40];
  assign d_o_t0[41] = _234_ | in_t0[41];
  assign d_o_t0[42] = _236_ | in_t0[42];
  assign d_o_t0[43] = _238_ | in_t0[43];
  assign d_o_t0[44] = _240_ | in_t0[44];
  assign d_o_t0[45] = _242_ | in_t0[45];
  assign d_o_t0[46] = _244_ | in_t0[46];
  assign d_o_t0[47] = _246_ | in_t0[47];
  assign d_o_t0[48] = _248_ | in_t0[48];
  assign d_o_t0[49] = _250_ | in_t0[49];
  assign d_o_t0[50] = _252_ | in_t0[50];
  assign d_o_t0[51] = _254_ | in_t0[51];
  assign d_o_t0[52] = _256_ | in_t0[52];
  assign d_o_t0[53] = _258_ | in_t0[53];
  assign d_o_t0[54] = _260_ | in_t0[54];
  assign d_o_t0[55] = _262_ | in_t0[55];
  assign d_o_t0[56] = _264_ | in_t0[56];
  assign _151_ = syndrome_o == 7'h07;
  assign _153_ = syndrome_o == 7'h0b;
  assign _155_ = syndrome_o == 7'h13;
  assign _157_ = syndrome_o == 7'h23;
  assign _159_ = syndrome_o == 7'h43;
  assign _161_ = syndrome_o == 7'h0d;
  assign _163_ = syndrome_o == 7'h15;
  assign _165_ = syndrome_o == 7'h25;
  assign _167_ = syndrome_o == 7'h45;
  assign _169_ = syndrome_o == 7'h19;
  assign _171_ = syndrome_o == 7'h29;
  assign _173_ = syndrome_o == 7'h49;
  assign _175_ = syndrome_o == 7'h31;
  assign _177_ = syndrome_o == 7'h51;
  assign _179_ = syndrome_o == 7'h61;
  assign _181_ = syndrome_o == 7'h0e;
  assign _183_ = syndrome_o == 7'h16;
  assign _185_ = syndrome_o == 7'h26;
  assign _187_ = syndrome_o == 7'h46;
  assign _189_ = syndrome_o == 7'h1a;
  assign _191_ = syndrome_o == 7'h2a;
  assign _193_ = syndrome_o == 7'h4a;
  assign _195_ = syndrome_o == 7'h32;
  assign _197_ = syndrome_o == 7'h52;
  assign _199_ = syndrome_o == 7'h62;
  assign _201_ = syndrome_o == 7'h1c;
  assign _203_ = syndrome_o == 7'h2c;
  assign _205_ = syndrome_o == 7'h4c;
  assign _207_ = syndrome_o == 7'h34;
  assign _209_ = syndrome_o == 7'h54;
  assign _211_ = syndrome_o == 7'h64;
  assign _213_ = syndrome_o == 7'h38;
  assign _215_ = syndrome_o == 7'h58;
  assign _217_ = syndrome_o == 7'h68;
  assign _219_ = syndrome_o == 7'h70;
  assign _221_ = syndrome_o == 7'h1f;
  assign _223_ = syndrome_o == 7'h2f;
  assign _225_ = syndrome_o == 7'h4f;
  assign _227_ = syndrome_o == 7'h37;
  assign _229_ = syndrome_o == 7'h57;
  assign _231_ = syndrome_o == 7'h67;
  assign _233_ = syndrome_o == 7'h3b;
  assign _235_ = syndrome_o == 7'h5b;
  assign _237_ = syndrome_o == 7'h6b;
  assign _239_ = syndrome_o == 7'h73;
  assign _241_ = syndrome_o == 7'h3d;
  assign _243_ = syndrome_o == 7'h5d;
  assign _245_ = syndrome_o == 7'h6d;
  assign _247_ = syndrome_o == 7'h75;
  assign _249_ = syndrome_o == 7'h79;
  assign _251_ = syndrome_o == 7'h3e;
  assign _253_ = syndrome_o == 7'h5e;
  assign _255_ = syndrome_o == 7'h6e;
  assign _257_ = syndrome_o == 7'h76;
  assign _259_ = syndrome_o == 7'h7a;
  assign _261_ = syndrome_o == 7'h7c;
  assign _263_ = syndrome_o == 7'h7f;
  assign _265_ = ~ single_error;
  assign _266_ = | syndrome_o;
  assign syndrome_o[0] = ^ _000_;
  assign syndrome_o[1] = ^ _002_;
  assign syndrome_o[2] = ^ _004_;
  assign syndrome_o[3] = ^ _006_;
  assign syndrome_o[4] = ^ _008_;
  assign syndrome_o[5] = ^ _010_;
  assign syndrome_o[6] = ^ _012_;
  assign single_error = ^ syndrome_o;
  assign d_o[0] = _151_ ^ in[0];
  assign d_o[1] = _153_ ^ in[1];
  assign d_o[2] = _155_ ^ in[2];
  assign d_o[3] = _157_ ^ in[3];
  assign d_o[4] = _159_ ^ in[4];
  assign d_o[5] = _161_ ^ in[5];
  assign d_o[6] = _163_ ^ in[6];
  assign d_o[7] = _165_ ^ in[7];
  assign d_o[8] = _167_ ^ in[8];
  assign d_o[9] = _169_ ^ in[9];
  assign d_o[10] = _171_ ^ in[10];
  assign d_o[11] = _173_ ^ in[11];
  assign d_o[12] = _175_ ^ in[12];
  assign d_o[13] = _177_ ^ in[13];
  assign d_o[14] = _179_ ^ in[14];
  assign d_o[15] = _181_ ^ in[15];
  assign d_o[16] = _183_ ^ in[16];
  assign d_o[17] = _185_ ^ in[17];
  assign d_o[18] = _187_ ^ in[18];
  assign d_o[19] = _189_ ^ in[19];
  assign d_o[20] = _191_ ^ in[20];
  assign d_o[21] = _193_ ^ in[21];
  assign d_o[22] = _195_ ^ in[22];
  assign d_o[23] = _197_ ^ in[23];
  assign d_o[24] = _199_ ^ in[24];
  assign d_o[25] = _201_ ^ in[25];
  assign d_o[26] = _203_ ^ in[26];
  assign d_o[27] = _205_ ^ in[27];
  assign d_o[28] = _207_ ^ in[28];
  assign d_o[29] = _209_ ^ in[29];
  assign d_o[30] = _211_ ^ in[30];
  assign d_o[31] = _213_ ^ in[31];
  assign d_o[32] = _215_ ^ in[32];
  assign d_o[33] = _217_ ^ in[33];
  assign d_o[34] = _219_ ^ in[34];
  assign d_o[35] = _221_ ^ in[35];
  assign d_o[36] = _223_ ^ in[36];
  assign d_o[37] = _225_ ^ in[37];
  assign d_o[38] = _227_ ^ in[38];
  assign d_o[39] = _229_ ^ in[39];
  assign d_o[40] = _231_ ^ in[40];
  assign d_o[41] = _233_ ^ in[41];
  assign d_o[42] = _235_ ^ in[42];
  assign d_o[43] = _237_ ^ in[43];
  assign d_o[44] = _239_ ^ in[44];
  assign d_o[45] = _241_ ^ in[45];
  assign d_o[46] = _243_ ^ in[46];
  assign d_o[47] = _245_ ^ in[47];
  assign d_o[48] = _247_ ^ in[48];
  assign d_o[49] = _249_ ^ in[49];
  assign d_o[50] = _251_ ^ in[50];
  assign d_o[51] = _253_ ^ in[51];
  assign d_o[52] = _255_ ^ in[52];
  assign d_o[53] = _257_ ^ in[53];
  assign d_o[54] = _259_ ^ in[54];
  assign d_o[55] = _261_ ^ in[55];
  assign d_o[56] = _263_ ^ in[56];
  assign err_o[0] = single_error;
  assign err_o_t0[0] = single_error_t0;
endmodule

module auxy_prim_secded_64_57_enc(in, out, in_t0, out_t0);
  wire [63:0] _00_;
  wire [63:0] _01_;
  wire [63:0] _02_;
  wire [63:0] _03_;
  wire [63:0] _04_;
  wire [63:0] _05_;
  wire [63:0] _06_;
  wire [63:0] _07_;
  wire [63:0] _08_;
  wire [63:0] _09_;
  wire [63:0] _10_;
  wire [63:0] _11_;
  wire [63:0] _12_;
  wire [63:0] _13_;
  wire [63:0] _14_;
  wire [63:0] _15_;
  wire [63:0] _16_;
  wire [63:0] _17_;
  wire [63:0] _18_;
  wire [63:0] _19_;
  wire [63:0] _20_;
  wire [63:0] _21_;
  wire [63:0] _22_;
  wire [63:0] _23_;
  wire [63:0] _24_;
  wire [63:0] _25_;
  wire [63:0] _26_;
  wire [63:0] _27_;
  wire [63:0] _28_;
  wire [63:0] _29_;
  wire [63:0] _30_;
  wire [63:0] _31_;
  wire [63:0] _32_;
  wire [63:0] _33_;
  wire [63:0] _34_;
  wire [63:0] _35_;
  wire [63:0] _36_;
  wire [63:0] _37_;
  wire [63:0] _38_;
  wire [63:0] _39_;
  wire [63:0] _40_;
  wire [63:0] _41_;
  input [56:0] in;
  wire [56:0] in;
  input [56:0] in_t0;
  wire [56:0] in_t0;
  output [63:0] out;
  wire [63:0] out;
  output [63:0] out_t0;
  wire [63:0] out_t0;
  assign _00_ = { 7'h00, in } & 64'h0103fff800007fff;
  assign _02_ = { 6'h00, out[57], in } & 64'h017c1ff801ff801f;
  assign _04_ = { 5'h00, out[58:57], in } & 64'h01bde1f87e0781e1;
  assign _06_ = { 4'h0, out[59:57], in } & 64'h01deee3b8e388e22;
  assign _08_ = { 3'h0, out[60:57], in } & 64'h01ef76cdb2c93244;
  assign _10_ = { 2'h0, out[61:57], in } & 64'h01f7bb56d5525488;
  assign _12_ = { 1'h0, out[62:57], in } & 64'h01fbdda769a46910;
  assign _14_ = { 7'h00, in_t0 } & 64'h0103fff800007fff;
  assign _17_ = { 6'h00, out_t0[57], in_t0 } & 64'h017c1ff801ff801f;
  assign _20_ = { 5'h00, out_t0[58:57], in_t0 } & 64'h01bde1f87e0781e1;
  assign _23_ = { 4'h0, out_t0[59:57], in_t0 } & 64'h01deee3b8e388e22;
  assign _26_ = { 3'h0, out_t0[60:57], in_t0 } & 64'h01ef76cdb2c93244;
  assign _29_ = { 2'h0, out_t0[61:57], in_t0 } & 64'h01f7bb56d5525488;
  assign _32_ = { 1'h0, out_t0[62:57], in_t0 } & 64'h01fbdda769a46910;
  assign _15_ = 64'h0000000000000000 & { 7'h00, in };
  assign _18_ = 64'h0000000000000000 & { 6'h00, out[57], in };
  assign _21_ = 64'h0000000000000000 & { 5'h00, out[58:57], in };
  assign _24_ = 64'h0000000000000000 & { 4'h0, out[59:57], in };
  assign _27_ = 64'h0000000000000000 & { 3'h0, out[60:57], in };
  assign _30_ = 64'h0000000000000000 & { 2'h0, out[61:57], in };
  assign _33_ = 64'h0000000000000000 & { 1'h0, out[62:57], in };
  assign _16_ = { 7'h00, in_t0 } & 64'h0000000000000000;
  assign _19_ = { 6'h00, out_t0[57], in_t0 } & 64'h0000000000000000;
  assign _22_ = { 5'h00, out_t0[58:57], in_t0 } & 64'h0000000000000000;
  assign _25_ = { 4'h0, out_t0[59:57], in_t0 } & 64'h0000000000000000;
  assign _28_ = { 3'h0, out_t0[60:57], in_t0 } & 64'h0000000000000000;
  assign _31_ = { 2'h0, out_t0[61:57], in_t0 } & 64'h0000000000000000;
  assign _34_ = { 1'h0, out_t0[62:57], in_t0 } & 64'h0000000000000000;
  assign _35_ = _14_ | _15_;
  assign _36_ = _17_ | _18_;
  assign _37_ = _20_ | _21_;
  assign _38_ = _23_ | _24_;
  assign _39_ = _26_ | _27_;
  assign _40_ = _29_ | _30_;
  assign _41_ = _32_ | _33_;
  assign _01_ = _35_ | _16_;
  assign _03_ = _36_ | _19_;
  assign _05_ = _37_ | _22_;
  assign _07_ = _38_ | _25_;
  assign _09_ = _39_ | _28_;
  assign _11_ = _40_ | _31_;
  assign _13_ = _41_ | _34_;
  assign out_t0[57] = | _01_;
  assign out_t0[58] = | _03_;
  assign out_t0[59] = | _05_;
  assign out_t0[60] = | _07_;
  assign out_t0[61] = | _09_;
  assign out_t0[62] = | _11_;
  assign out_t0[63] = | _13_;
  assign out[57] = ^ _00_;
  assign out[58] = ^ _02_;
  assign out[59] = ^ _04_;
  assign out[60] = ^ _06_;
  assign out[61] = ^ _08_;
  assign out[62] = ^ _10_;
  assign out[63] = ^ _12_;
  assign out[56:0] = in;
  assign out_t0[56:0] = in_t0;
endmodule

module auxy_rv_core_ibex_mem_top(clk_i, rst_ni, clk_esc_i, rst_esc_ni, test_en_i, ram_cfg_i, hart_id_i, boot_addr_i, instr_mem_req_o, instr_mem_gnt_i, instr_mem_addr_o, instr_mem_wdata_o, instr_mem_strb_o, instr_mem_we_o, instr_mem_rdata_i, data_mem_req_o, data_mem_gnt_i, data_mem_addr_o, data_mem_wdata_o, data_mem_strb_o, data_mem_we_o
, data_mem_rdata_i, irq_software_i, irq_timer_i, irq_external_i, esc_tx_i, esc_rx_o, debug_req_i, crash_dump_o, lc_cpu_en_i, core_sleep_o, boot_addr_i_t0, test_en_i_t0, esc_rx_o_t0, esc_tx_i_t0, debug_req_i_t0, hart_id_i_t0, irq_external_i_t0, irq_software_i_t0, irq_timer_i_t0, crash_dump_o_t0, core_sleep_o_t0
, ram_cfg_i_t0, clk_esc_i_t0, lc_cpu_en_i_t0, rst_esc_ni_t0, data_mem_addr_o_t0, data_mem_gnt_i_t0, data_mem_rdata_i_t0, data_mem_req_o_t0, data_mem_strb_o_t0, data_mem_wdata_o_t0, data_mem_we_o_t0, instr_mem_addr_o_t0, instr_mem_gnt_i_t0, instr_mem_rdata_i_t0, instr_mem_req_o_t0, instr_mem_strb_o_t0, instr_mem_wdata_o_t0, instr_mem_we_o_t0);
  wire _00_;
  wire _01_;
  wire _02_;
  wire _03_;
  wire _04_;
  wire _05_;
  wire _06_;
  wire _07_;
  wire _08_;
  wire _09_;
  input [31:0] boot_addr_i /* verilator public */;
  wire [31:0] boot_addr_i;
  input [31:0] boot_addr_i_t0 /* verilator public */;
  wire [31:0] boot_addr_i_t0;
  input clk_esc_i /* verilator public */;
  wire clk_esc_i;
  input clk_esc_i_t0 /* verilator public */;
  wire clk_esc_i_t0;
  input clk_i /* verilator public */;
  wire clk_i;
  output core_sleep_o;
  wire core_sleep_o;
  output core_sleep_o_t0;
  wire core_sleep_o_t0;
  output [127:0] crash_dump_o;
  wire [127:0] crash_dump_o;
  output [127:0] crash_dump_o_t0;
  wire [127:0] crash_dump_o_t0;
  output [17:0] data_mem_addr_o;
  wire [17:0] data_mem_addr_o;
  output [17:0] data_mem_addr_o_t0;
  wire [17:0] data_mem_addr_o_t0;
  input data_mem_gnt_i /* verilator public */;
  wire data_mem_gnt_i;
  input data_mem_gnt_i_t0 /* verilator public */;
  wire data_mem_gnt_i_t0;
  input [31:0] data_mem_rdata_i /* verilator public */;
  wire [31:0] data_mem_rdata_i;
  input [31:0] data_mem_rdata_i_t0 /* verilator public */;
  wire [31:0] data_mem_rdata_i_t0;
  output data_mem_req_o;
  wire data_mem_req_o;
  output data_mem_req_o_t0;
  wire data_mem_req_o_t0;
  output [31:0] data_mem_strb_o;
  wire [31:0] data_mem_strb_o;
  output [31:0] data_mem_strb_o_t0;
  wire [31:0] data_mem_strb_o_t0;
  output [31:0] data_mem_wdata_o;
  wire [31:0] data_mem_wdata_o;
  output [31:0] data_mem_wdata_o_t0;
  wire [31:0] data_mem_wdata_o_t0;
  output data_mem_we_o;
  wire data_mem_we_o;
  output data_mem_we_o_t0;
  wire data_mem_we_o_t0;
  wire data_rvalid_d;
  wire data_rvalid_d_t0;
  reg data_rvalid_q;
  reg data_rvalid_q_t0;
  input debug_req_i /* verilator public */;
  wire debug_req_i;
  input debug_req_i_t0 /* verilator public */;
  wire debug_req_i_t0;
  output [1:0] esc_rx_o;
  wire [1:0] esc_rx_o;
  output [1:0] esc_rx_o_t0;
  wire [1:0] esc_rx_o_t0;
  input [1:0] esc_tx_i /* verilator public */;
  wire [1:0] esc_tx_i;
  input [1:0] esc_tx_i_t0 /* verilator public */;
  wire [1:0] esc_tx_i_t0;
  input [31:0] hart_id_i /* verilator public */;
  wire [31:0] hart_id_i;
  input [31:0] hart_id_i_t0 /* verilator public */;
  wire [31:0] hart_id_i_t0;
  output [17:0] instr_mem_addr_o;
  wire [17:0] instr_mem_addr_o;
  output [17:0] instr_mem_addr_o_t0;
  wire [17:0] instr_mem_addr_o_t0;
  input instr_mem_gnt_i /* verilator public */;
  wire instr_mem_gnt_i;
  input instr_mem_gnt_i_t0 /* verilator public */;
  wire instr_mem_gnt_i_t0;
  input [31:0] instr_mem_rdata_i /* verilator public */;
  wire [31:0] instr_mem_rdata_i;
  input [31:0] instr_mem_rdata_i_t0 /* verilator public */;
  wire [31:0] instr_mem_rdata_i_t0;
  output instr_mem_req_o;
  wire instr_mem_req_o;
  output instr_mem_req_o_t0;
  wire instr_mem_req_o_t0;
  output [31:0] instr_mem_strb_o;
  wire [31:0] instr_mem_strb_o;
  output [31:0] instr_mem_strb_o_t0;
  wire [31:0] instr_mem_strb_o_t0;
  output [31:0] instr_mem_wdata_o;
  wire [31:0] instr_mem_wdata_o;
  output [31:0] instr_mem_wdata_o_t0;
  wire [31:0] instr_mem_wdata_o_t0;
  output instr_mem_we_o;
  wire instr_mem_we_o;
  output instr_mem_we_o_t0;
  wire instr_mem_we_o_t0;
  wire instr_rvalid_d;
  wire instr_rvalid_d_t0;
  reg instr_rvalid_q;
  reg instr_rvalid_q_t0;
  input irq_external_i /* verilator public */;
  wire irq_external_i;
  input irq_external_i_t0 /* verilator public */;
  wire irq_external_i_t0;
  input irq_software_i /* verilator public */;
  wire irq_software_i;
  input irq_software_i_t0 /* verilator public */;
  wire irq_software_i_t0;
  input irq_timer_i /* verilator public */;
  wire irq_timer_i;
  input irq_timer_i_t0 /* verilator public */;
  wire irq_timer_i_t0;
  input [3:0] lc_cpu_en_i /* verilator public */;
  wire [3:0] lc_cpu_en_i;
  input [3:0] lc_cpu_en_i_t0 /* verilator public */;
  wire [3:0] lc_cpu_en_i_t0;
  input [9:0] ram_cfg_i /* verilator public */;
  wire [9:0] ram_cfg_i;
  input [9:0] ram_cfg_i_t0 /* verilator public */;
  wire [9:0] ram_cfg_i_t0;
  input rst_esc_ni /* verilator public */;
  wire rst_esc_ni;
  input rst_esc_ni_t0 /* verilator public */;
  wire rst_esc_ni_t0;
  input rst_ni /* verilator public */;
  wire rst_ni;
  input test_en_i /* verilator public */;
  wire test_en_i;
  input test_en_i_t0 /* verilator public */;
  wire test_en_i_t0;
  wire [106:0] tl_d_fromibex;
  wire [106:0] tl_d_fromibex_t0;
  wire [65:0] tl_d_toibex;
  wire [65:0] tl_d_toibex_t0;
  wire [106:0] tl_i_fromibex;
  wire [106:0] tl_i_fromibex_t0;
  wire [65:0] tl_i_toibex;
  wire [65:0] tl_i_toibex_t0;
  assign instr_rvalid_d = instr_mem_req_o & _08_;
  assign data_rvalid_d = data_mem_req_o & _09_;
  assign _00_ = instr_mem_req_o_t0 & _08_;
  assign _03_ = data_mem_req_o_t0 & _09_;
  assign _01_ = instr_mem_we_o_t0 & instr_mem_req_o;
  assign _04_ = data_mem_we_o_t0 & data_mem_req_o;
  assign _02_ = instr_mem_req_o_t0 & instr_mem_we_o_t0;
  assign _05_ = data_mem_req_o_t0 & data_mem_we_o_t0;
  assign _06_ = _00_ | _01_;
  assign _07_ = _03_ | _04_;
  assign instr_rvalid_d_t0 = _06_ | _02_;
  assign data_rvalid_d_t0 = _07_ | _05_;
  always_ff @(posedge clk_i)
    if (!rst_ni) instr_rvalid_q <= 1'h0;
    else instr_rvalid_q <= instr_rvalid_d;
  always_ff @(posedge clk_i)
    if (!rst_ni) data_rvalid_q <= 1'h0;
    else data_rvalid_q <= data_rvalid_d;
  always_ff @(posedge clk_i)
    if (!rst_ni) instr_rvalid_q_t0 <= 1'h0;
    else instr_rvalid_q_t0 <= instr_rvalid_d_t0;
  always_ff @(posedge clk_i)
    if (!rst_ni) data_rvalid_q_t0 <= 1'h0;
    else data_rvalid_q_t0 <= data_rvalid_d_t0;
  assign _08_ = ~ instr_mem_we_o;
  assign _09_ = ~ data_mem_we_o;
  paramodb14a8c3636c7c0bb82862600beccd3d8da4d4a94auxy_noerr_tlul_adapter_sram  i_data_tlul_adapter_sram (
    .addr_o(data_mem_addr_o),
    .addr_o_t0(data_mem_addr_o_t0),
    .clk_i(clk_i),
    .en_ifetch_i(3'h5),
    .en_ifetch_i_t0(3'h0),
    .gnt_i(data_mem_gnt_i),
    .gnt_i_t0(data_mem_gnt_i_t0),
    .rdata_i(data_mem_rdata_i),
    .rdata_i_t0(data_mem_rdata_i_t0),
    .req_o(data_mem_req_o),
    .req_o_t0(data_mem_req_o_t0),
    .rerror_i(2'h0),
    .rerror_i_t0(2'h0),
    .rst_ni(rst_ni),
    .rvalid_i(data_rvalid_q),
    .rvalid_i_t0(data_rvalid_q_t0),
    .tl_i(tl_d_fromibex),
    .tl_i_t0(tl_d_fromibex_t0),
    .tl_o(tl_d_toibex),
    .tl_o_t0(tl_d_toibex_t0),
    .wdata_o(data_mem_wdata_o),
    .wdata_o_t0(data_mem_wdata_o_t0),
    .we_o(data_mem_we_o),
    .we_o_t0(data_mem_we_o_t0),
    .wmask_o(data_mem_strb_o),
    .wmask_o_t0(data_mem_strb_o_t0)
  );
  paramodb14a8c3636c7c0bb82862600beccd3d8da4d4a94auxy_noerr_tlul_adapter_sram  i_instr_tlul_adapter_sram (
    .addr_o(instr_mem_addr_o),
    .addr_o_t0(instr_mem_addr_o_t0),
    .clk_i(clk_i),
    .en_ifetch_i(3'h5),
    .en_ifetch_i_t0(3'h0),
    .gnt_i(instr_mem_gnt_i),
    .gnt_i_t0(instr_mem_gnt_i_t0),
    .rdata_i(instr_mem_rdata_i),
    .rdata_i_t0(instr_mem_rdata_i_t0),
    .req_o(instr_mem_req_o),
    .req_o_t0(instr_mem_req_o_t0),
    .rerror_i(2'h0),
    .rerror_i_t0(2'h0),
    .rst_ni(rst_ni),
    .rvalid_i(instr_rvalid_q),
    .rvalid_i_t0(instr_rvalid_q_t0),
    .tl_i(tl_i_fromibex),
    .tl_i_t0(tl_i_fromibex_t0),
    .tl_o(tl_i_toibex),
    .tl_o_t0(tl_i_toibex_t0),
    .wdata_o(instr_mem_wdata_o),
    .wdata_o_t0(instr_mem_wdata_o_t0),
    .we_o(instr_mem_we_o),
    .we_o_t0(instr_mem_we_o_t0),
    .wmask_o(instr_mem_strb_o),
    .wmask_o_t0(instr_mem_strb_o_t0)
  );
  auxy_noerr_rv_core_ibex i_rv_core_ibex (
    .boot_addr_i(boot_addr_i),
    .boot_addr_i_t0(boot_addr_i_t0),
    .clk_esc_i(clk_esc_i),
    .clk_esc_i_t0(clk_esc_i_t0),
    .clk_i(clk_i),
    .core_sleep_o(core_sleep_o),
    .core_sleep_o_t0(core_sleep_o_t0),
    .crash_dump_o(crash_dump_o),
    .crash_dump_o_t0(crash_dump_o_t0),
    .debug_req_i(debug_req_i),
    .debug_req_i_t0(debug_req_i_t0),
    .esc_rx_o(esc_rx_o),
    .esc_rx_o_t0(esc_rx_o_t0),
    .esc_tx_i(esc_tx_i),
    .esc_tx_i_t0(esc_tx_i_t0),
    .hart_id_i(hart_id_i),
    .hart_id_i_t0(hart_id_i_t0),
    .irq_external_i(irq_external_i),
    .irq_external_i_t0(irq_external_i_t0),
    .irq_software_i(irq_software_i),
    .irq_software_i_t0(irq_software_i_t0),
    .irq_timer_i(irq_timer_i),
    .irq_timer_i_t0(irq_timer_i_t0),
    .lc_cpu_en_i(lc_cpu_en_i),
    .lc_cpu_en_i_t0(lc_cpu_en_i_t0),
    .ram_cfg_i(ram_cfg_i),
    .ram_cfg_i_t0(ram_cfg_i_t0),
    .rst_esc_ni(rst_esc_ni),
    .rst_esc_ni_t0(rst_esc_ni_t0),
    .rst_ni(rst_ni),
    .test_en_i(test_en_i),
    .test_en_i_t0(test_en_i_t0),
    .tl_d_i(tl_d_toibex),
    .tl_d_i_t0(tl_d_toibex_t0),
    .tl_d_o(tl_d_fromibex),
    .tl_d_o_t0(tl_d_fromibex_t0),
    .tl_i_i(tl_i_toibex),
    .tl_i_i_t0(tl_i_toibex_t0),
    .tl_i_o(tl_i_fromibex),
    .tl_i_o_t0(tl_i_fromibex_t0)
  );
endmodule

module auxy_tlul_cmd_intg_gen(tl_i, tl_o, tl_i_t0, tl_o_t0);
  input [106:0] tl_i;
  wire [106:0] tl_i;
  input [106:0] tl_i_t0;
  wire [106:0] tl_i_t0;
  output [106:0] tl_o;
  wire [106:0] tl_o;
  output [106:0] tl_o_t0;
  wire [106:0] tl_o_t0;
  wire [56:0] unused_cmd_payload;
  wire [56:0] unused_cmd_payload_t0;
  auxy_prim_secded_64_57_enc u_cmd_gen (
    .in({ 16'h0000, tl_i[16:15], tl_i[89:58], tl_i[105:103], tl_i[57:54] }),
    .in_t0({ 16'h0000, tl_i_t0[16:15], tl_i_t0[89:58], tl_i_t0[105:103], tl_i_t0[57:54] }),
    .out({ tl_o[14:8], unused_cmd_payload }),
    .out_t0({ tl_o_t0[14:8], unused_cmd_payload_t0 })
  );
  assign { tl_o[106:15], tl_o[7:0] } = { tl_i[106:15], tl_i[7:0] };
  assign { tl_o_t0[106:15], tl_o_t0[7:0] } = { tl_i_t0[106:15], tl_i_t0[7:0] };
endmodule





module auxy_tlul_rsp_intg_chk(tl_i, err_o, err_o_t0, tl_i_t0);
  wire [1:0] _00_;
  wire _01_;
  wire _02_;
  wire _03_;
  wire _04_;
  wire _05_;
  wire [1:0] _06_;
  wire _07_;
  wire _08_;
  wire _09_;
  wire [1:0] err;
  output err_o;
  wire err_o;
  output err_o_t0;
  wire err_o_t0;
  wire [1:0] err_t0;
  input [65:0] tl_i;
  wire [65:0] tl_i;
  input [65:0] tl_i_t0;
  wire [65:0] tl_i_t0;
  assign err_o = tl_i[65] & _08_;
  assign _03_ = tl_i_t0[65] & _08_;
  assign _04_ = _09_ & tl_i[65];
  assign _05_ = tl_i_t0[65] & _09_;
  assign _07_ = _03_ | _04_;
  assign err_o_t0 = _07_ | _05_;
  assign _01_ = | err_t0;
  assign _00_ = ~ err_t0;
  assign _06_ = err & _00_;
  assign _02_ = ! _06_;
  assign _09_ = _02_ & _01_;
  assign _08_ = | err;
  auxy_prim_secded_64_57_dec u_chk (
    .err_o(err),
    .err_o_t0(err_t0),
    .in({ tl_i[15:9], 51'h0000000000000, tl_i[64:62], tl_i[58:57], tl_i[1] }),
    .in_t0({ tl_i_t0[15:9], 51'h0000000000000, tl_i_t0[64:62], tl_i_t0[58:57], tl_i_t0[1] })
  );
endmodule

